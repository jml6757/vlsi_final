//
// Verilog description for cell filter, 
// Fri Dec 12 16:11:30 2014
//
// LeonardoSpectrum Level 3, 2008b.3 
//


module filter ( T00, T01, T02, T10, T11, T12, T20, T21, T22, CLOCK, I_VALID, 
                RESET, THRESHOLD, READY, O_VALID, EDGE, DIRECTION ) ;

    input [7:0]T00 ;
    input [7:0]T01 ;
    input [7:0]T02 ;
    input [7:0]T10 ;
    input [7:0]T11 ;
    input [7:0]T12 ;
    input [7:0]T20 ;
    input [7:0]T21 ;
    input [7:0]T22 ;
    input CLOCK ;
    input I_VALID ;
    input RESET ;
    input [10:0]THRESHOLD ;
    output READY ;
    output O_VALID ;
    output EDGE ;
    output [2:0]DIRECTION ;

    wire nx1586, fsm_inst_state_3, fsm_inst_state_2, fsm_inst_state_0, nx8, nx12, 
         nx18, nx56, nx70, nx78, nx88, nx94, nx104, nx110, nx120, nx126, nx128, 
         nx140, nx150, nx158, nx166, nx174, nx182, nx192, nx220, nx234, nx242, 
         nx252, nx258, nx268, nx274, nx284, nx290, nx292, nx304, nx314, nx322, 
         nx330, nx338, nx346, nx356, nx360, nx368, nx374, nx380, nx392, nx398, 
         nx400, nx408, nx410, nx412, nx420, nx422, nx424, nx432, nx434, nx436, 
         nx444, nx446, nx448, nx456, nx458, nx460, nx472, nx480, nx482, nx484, 
         nx510, nx518, nx526, nx534, nx542, nx544, nx608, nx616, nx624, nx632, 
         nx640, nx646, nx678, nx692, nx700, nx710, nx716, nx726, nx732, nx742, 
         nx748, nx750, nx762, nx772, nx780, nx788, nx796, nx804, nx814, nx842, 
         nx856, nx864, nx874, nx880, nx890, nx896, nx906, nx912, nx914, nx926, 
         nx936, nx944, nx952, nx960, nx968, nx978, nx990, nx996, nx1002, nx1014, 
         nx1020, nx1022, nx1030, nx1032, nx1034, nx1042, nx1044, nx1046, nx1054, 
         nx1056, nx1058, nx1066, nx1068, nx1070, nx1078, nx1080, nx1082, nx1094, 
         nx1102, nx1104, nx1106, nx1132, nx1140, nx1148, nx1156, nx1164, nx1166, 
         nx1230, nx1238, nx1246, nx1254, nx1262, nx1268, nx1278, nx1284, nx1288, 
         nx1290, nx1296, nx1314, nx1326, nx1330, nx1336, nx1340, nx1342, nx1348, 
         nx1366, nx1378, nx1382, nx1388, nx1392, nx1394, nx1400, nx1418, nx1430, 
         nx1434, nx1440, nx1444, nx1446, nx1452, nx1470, nx1482, nx1486, nx1492, 
         nx1498, nx1504, nx1516, nx1534, nx1550, nx1566, nx1582, nx1598, nx1640, 
         nx1654, nx1662, nx1672, nx1678, nx1688, nx1694, nx1704, nx1710, nx1712, 
         nx1724, nx1734, nx1742, nx1750, nx1758, nx1766, nx1776, nx1804, nx1818, 
         nx1826, nx1836, nx1842, nx1852, nx1858, nx1868, nx1874, nx1876, nx1888, 
         nx1898, nx1906, nx1914, nx1922, nx1930, nx1940, nx1952, nx1958, nx1964, 
         nx1976, nx1982, nx1984, nx1992, nx1994, nx1996, nx2004, nx2006, nx2008, 
         nx2016, nx2018, nx2020, nx2028, nx2030, nx2032, nx2040, nx2042, nx2044, 
         nx2056, nx2064, nx2066, nx2068, nx2094, nx2102, nx2110, nx2118, nx2126, 
         nx2128, nx2192, nx2200, nx2208, nx2216, nx2224, nx2230, nx2262, nx2276, 
         nx2284, nx2294, nx2300, nx2310, nx2316, nx2326, nx2332, nx2334, nx2346, 
         nx2356, nx2364, nx2372, nx2380, nx2388, nx2398, nx2426, nx2440, nx2448, 
         nx2458, nx2464, nx2474, nx2480, nx2490, nx2496, nx2498, nx2510, nx2520, 
         nx2528, nx2536, nx2544, nx2552, nx2562, nx2574, nx2580, nx2586, nx2598, 
         nx2604, nx2606, nx2614, nx2616, nx2618, nx2626, nx2628, nx2630, nx2638, 
         nx2640, nx2642, nx2650, nx2652, nx2654, nx2662, nx2664, nx2666, nx2678, 
         nx2686, nx2688, nx2690, nx2716, nx2724, nx2732, nx2740, nx2748, nx2750, 
         nx2814, nx2822, nx2830, nx2838, nx2846, nx2852, nx2862, nx2868, nx2874, 
         nx2880, nx2884, nx2898, nx2910, nx2914, nx2920, nx2926, nx2932, nx2936, 
         nx2950, nx2962, nx2966, nx2972, nx2978, nx2984, nx2988, nx3002, nx3014, 
         nx3018, nx3024, nx3030, nx3036, nx3040, nx3054, nx3066, nx3070, nx3076, 
         nx3082, nx3088, nx3100, nx3118, nx3134, nx3150, nx3166, nx3182, nx3208, 
         nx3216, nx3244, nx3252, nx3280, nx3288, nx3316, nx3324, nx3352, nx3360, 
         nx3370, nx3378, nx3382, nx3398, nx3414, nx3430, nx3446, nx3462, nx3466, 
         nx3472, nx3478, nx3486, nx3490, nx3518, nx3520, nx3528, nx3530, nx3546, 
         nx3574, nx3576, nx3584, nx3586, nx3602, nx3630, nx3632, nx3640, nx3642, 
         nx3658, nx3694, nx3698, nx3702, nx3710, nx3718, nx3726, nx3734, nx3746, 
         nx3754, nx3758, nx3766, nx3774, nx3778, nx3782, nx3786, nx3790, nx3794, 
         nx3798, nx3800, nx3802, nx3820, nx3828, nx3836, nx3844, nx3852, nx3860, 
         nx3868, nx3876, nx3884, nx3904, nx1683, nx1691, nx1695, nx1699, nx1703, 
         nx1709, nx1711, nx1713, nx1715, nx1717, nx1719, nx1721, nx1723, nx1729, 
         nx1731, nx1735, nx1737, nx1741, nx1743, nx1747, nx1749, nx1753, nx1755, 
         nx1761, nx1767, nx1773, nx1779, nx1781, nx1783, nx1789, nx1791, nx1797, 
         nx1799, nx1805, nx1807, nx1813, nx1815, nx1817, nx1819, nx1827, nx1829, 
         nx1833, nx1839, nx1841, nx1847, nx1853, nx1855, nx1861, nx1869, nx1875, 
         nx1877, nx1885, nx1889, nx1891, nx1893, nx1901, nx1907, nx1909, nx1917, 
         nx1921, nx1923, nx1925, nx1933, nx1937, nx1943, nx1949, nx1951, nx1957, 
         nx1969, nx1971, nx1975, nx1977, nx1981, nx1983, nx1987, nx1991, nx1995, 
         nx2001, nx2007, nx2011, nx2013, nx2017, nx2023, nx2027, nx2029, nx2033, 
         nx2039, nx2043, nx2045, nx2049, nx2055, nx2059, nx2061, nx2065, nx2071, 
         nx2075, nx2077, nx2079, nx2081, nx2083, nx2085, nx2087, nx2089, nx2091, 
         nx2101, nx2103, nx2109, nx2111, nx2115, nx2123, nx2127, nx2131, nx2135, 
         nx2139, nx2141, nx2143, nx2145, nx2147, nx2149, nx2151, nx2153, nx2159, 
         nx2161, nx2165, nx2167, nx2171, nx2173, nx2177, nx2183, nx2189, nx2195, 
         nx2201, nx2203, nx2205, nx2211, nx2213, nx2219, nx2221, nx2227, nx2229, 
         nx2235, nx2241, nx2243, nx2249, nx2255, nx2257, nx2263, nx2271, nx2277, 
         nx2279, nx2287, nx2291, nx2293, nx2295, nx2303, nx2309, nx2311, nx2319, 
         nx2323, nx2325, nx2327, nx2335, nx2339, nx2345, nx2351, nx2353, nx2361, 
         nx2365, nx2367, nx2371, nx2373, nx2379, nx2381, nx2385, nx2387, nx2391, 
         nx2393, nx2399, nx2401, nx2403, nx2407, nx2409, nx2413, nx2415, nx2421, 
         nx2423, nx2425, nx2429, nx2431, nx2435, nx2437, nx2443, nx2445, nx2447, 
         nx2465, nx2475, nx2479, nx2483, nx2487, nx2491, nx2493, nx2495, nx2497, 
         nx2499, nx2501, nx2503, nx2505, nx2507, nx2513, nx2515, nx2519, nx2521, 
         nx2525, nx2527, nx2531, nx2533, nx2537, nx2539, nx2545, nx2551, nx2557, 
         nx2563, nx2565, nx2567, nx2573, nx2575, nx2579, nx2581, nx2587, nx2589, 
         nx2595, nx2597, nx2599, nx2601, nx2609, nx2611, nx2615, nx2621, nx2623, 
         nx2629, nx2635, nx2637, nx2641, nx2649, nx2655, nx2663, nx2667, nx2669, 
         nx2671, nx2679, nx2685, nx2693, nx2697, nx2699, nx2701, nx2709, nx2717, 
         nx2723, nx2725, nx2739, nx2741, nx2745, nx2747, nx2751, nx2753, nx2757, 
         nx2761, nx2769, nx2773, nx2777, nx2781, nx2787, nx2789, nx2791, nx2793, 
         nx2795, nx2797, nx2799, nx2805, nx2807, nx2811, nx2813, nx2817, nx2819, 
         nx2823, nx2825, nx2829, nx2831, nx2837, nx2843, nx2849, nx2855, nx2857, 
         nx2859, nx2865, nx2867, nx2873, nx2875, nx2879, nx2881, nx2887, nx2889, 
         nx2891, nx2893, nx2901, nx2903, nx2907, nx2913, nx2915, nx2919, nx2925, 
         nx2927, nx2933, nx2941, nx2945, nx2947, nx2955, nx2959, nx2961, nx2963, 
         nx2971, nx2977, nx2979, nx2985, nx2989, nx2991, nx2993, nx2999, nx3003, 
         nx3009, nx3015, nx3017, nx3031, nx3033, nx3037, nx3039, nx3043, nx3045, 
         nx3049, nx3053, nx3055, nx3059, nx3065, nx3071, nx3075, nx3081, nx3085, 
         nx3089, nx3091, nx3095, nx3101, nx3105, nx3107, nx3111, nx3117, nx3121, 
         nx3123, nx3127, nx3133, nx3137, nx3139, nx3143, nx3149, nx3153, nx3155, 
         nx3157, nx3163, nx3167, nx3169, nx3171, nx3173, nx3179, nx3183, nx3185, 
         nx3187, nx3189, nx3195, nx3199, nx3201, nx3203, nx3205, nx3211, nx3215, 
         nx3217, nx3219, nx3221, nx3225, nx3227, nx3231, nx3233, nx3239, nx3241, 
         nx3247, nx3249, nx3257, nx3261, nx3263, nx3267, nx3269, nx3271, nx3275, 
         nx3277, nx3279, nx3283, nx3285, nx3287, nx3291, nx3293, nx3295, nx3299, 
         nx3301, nx3307, nx3313, nx3319, nx3323, nx3327, nx3335, nx3357, nx3381, 
         nx3405, nx3407, nx3409, nx3429, nx3433, nx3435, nx3441, nx3461, nx3465, 
         nx3467, nx3473, nx3493, nx3497, nx3499, nx3505, nx3525, nx3537, nx3539, 
         nx3543, nx3547, nx3553, nx3555, nx3561, nx3563, nx3569, nx3571, nx3577, 
         nx3579, nx3587, nx3589, nx3595, nx3601, nx3607, nx3613, nx3619, nx3623, 
         nx3627, nx3631, nx3635, nx3641, nx3680, nx3686, nx3688, nx3690, nx3715, 
         nx3717, nx3719, nx3721, nx3727, nx3729, nx3731, nx3733, nx3735, nx3737, 
         nx3739, nx3741;
    wire [4:0] \$dummy ;




    fake_vcc ix1676 (.Y (nx360)) ;
    fake_gnd ix1587 (.Y (nx1586)) ;
    nor02ii ix3909 (.Y (DIRECTION[0]), .A0 (nx1683), .A1 (EDGE)) ;
    aoi221 ix1684 (.Y (nx1683), .A0 (nx3733), .A1 (nx3688), .B0 (nx3729), .B1 (
           nx3686), .C0 (nx3904)) ;
    mux21 ix2749 (.Y (nx2748), .A0 (nx2574), .A1 (nx1779), .S0 (nx2586)) ;
    nand02 ix1692 (.Y (nx1691), .A0 (T12[7]), .A1 (nx2388)) ;
    mux21 ix2389 (.Y (nx2388), .A0 (nx1695), .A1 (nx1721), .S0 (nx1723)) ;
    mux21 ix1696 (.Y (nx1695), .A0 (nx2284), .A1 (T02[6]), .S0 (nx1719)) ;
    mux21 ix2285 (.Y (nx2284), .A0 (nx1699), .A1 (nx1715), .S0 (nx1717)) ;
    mux21 ix1700 (.Y (nx1699), .A0 (nx2276), .A1 (T02[4]), .S0 (nx1713)) ;
    mux21 ix2277 (.Y (nx2276), .A0 (nx1703), .A1 (nx1709), .S0 (nx1711)) ;
    aoi32 ix1704 (.Y (nx1703), .A0 (T12[0]), .A1 (T02[1]), .A2 (nx2262), .B0 (
          T02[2]), .B1 (T12[1])) ;
    inv01 ix1710 (.Y (nx1709), .A (T02[3])) ;
    xnor2 ix1712 (.Y (nx1711), .A0 (T12[2]), .A1 (T02[3])) ;
    xnor2 ix1714 (.Y (nx1713), .A0 (T12[3]), .A1 (T02[4])) ;
    inv01 ix1716 (.Y (nx1715), .A (T02[5])) ;
    xnor2 ix1718 (.Y (nx1717), .A0 (T12[4]), .A1 (T02[5])) ;
    xnor2 ix1720 (.Y (nx1719), .A0 (T12[5]), .A1 (T02[6])) ;
    inv01 ix1722 (.Y (nx1721), .A (T02[7])) ;
    xnor2 ix1724 (.Y (nx1723), .A0 (T12[6]), .A1 (T02[7])) ;
    mux21 ix2381 (.Y (nx2380), .A0 (nx1729), .A1 (nx1731), .S0 (nx2294)) ;
    xnor2 ix1730 (.Y (nx1729), .A0 (nx1695), .A1 (nx1723)) ;
    mux21 ix1732 (.Y (nx1731), .A0 (nx2372), .A1 (nx2300), .S0 (nx1773)) ;
    mux21 ix2373 (.Y (nx2372), .A0 (nx1735), .A1 (nx1737), .S0 (nx2310)) ;
    xnor2 ix1736 (.Y (nx1735), .A0 (nx1699), .A1 (nx1717)) ;
    mux21 ix1738 (.Y (nx1737), .A0 (nx2364), .A1 (nx2316), .S0 (nx1767)) ;
    mux21 ix2365 (.Y (nx2364), .A0 (nx1741), .A1 (nx1743), .S0 (nx2326)) ;
    xnor2 ix1742 (.Y (nx1741), .A0 (nx1703), .A1 (nx1711)) ;
    aoi22 ix1744 (.Y (nx1743), .A0 (nx2332), .A1 (T22[2]), .B0 (nx2356), .B1 (
          nx2334)) ;
    nand02 ix1748 (.Y (nx1747), .A0 (T12[0]), .A1 (T02[1])) ;
    xnor2 ix1750 (.Y (nx1749), .A0 (T12[1]), .A1 (T02[2])) ;
    mux21 ix2357 (.Y (nx2356), .A0 (nx1753), .A1 (nx1755), .S0 (nx2346)) ;
    oai21 ix1754 (.Y (nx1753), .A0 (T02[1]), .A1 (T12[0]), .B0 (nx1747)) ;
    nand02 ix1756 (.Y (nx1755), .A0 (T22[0]), .A1 (T02[0])) ;
    xnor2 ix2347 (.Y (nx2346), .A0 (T22[1]), .A1 (nx1753)) ;
    xnor2 ix2335 (.Y (nx2334), .A0 (T22[2]), .A1 (nx1761)) ;
    xnor2 ix1762 (.Y (nx1761), .A0 (nx1747), .A1 (nx1749)) ;
    xnor2 ix2327 (.Y (nx2326), .A0 (T22[3]), .A1 (nx1741)) ;
    xnor2 ix2317 (.Y (nx2316), .A0 (nx2276), .A1 (nx1713)) ;
    xnor2 ix1768 (.Y (nx1767), .A0 (T22[4]), .A1 (nx2316)) ;
    xnor2 ix2311 (.Y (nx2310), .A0 (T22[5]), .A1 (nx1735)) ;
    xnor2 ix2301 (.Y (nx2300), .A0 (nx2284), .A1 (nx1719)) ;
    xnor2 ix1774 (.Y (nx1773), .A0 (T22[6]), .A1 (nx2300)) ;
    xnor2 ix2295 (.Y (nx2294), .A0 (T22[7]), .A1 (nx1729)) ;
    mux21 ix1780 (.Y (nx1779), .A0 (nx1781), .A1 (nx2740), .S0 (nx2606)) ;
    xnor2 ix1784 (.Y (nx1783), .A0 (T12[7]), .A1 (nx2388)) ;
    mux21 ix2741 (.Y (nx2740), .A0 (nx2614), .A1 (nx1789), .S0 (nx2618)) ;
    xnor2 ix2615 (.Y (nx2614), .A0 (nx1731), .A1 (nx2294)) ;
    mux21 ix1790 (.Y (nx1789), .A0 (nx1791), .A1 (nx2732), .S0 (nx2630)) ;
    mux21 ix2733 (.Y (nx2732), .A0 (nx2638), .A1 (nx1797), .S0 (nx2642)) ;
    xnor2 ix2639 (.Y (nx2638), .A0 (nx1737), .A1 (nx2310)) ;
    mux21 ix1798 (.Y (nx1797), .A0 (nx1799), .A1 (nx2724), .S0 (nx2654)) ;
    mux21 ix2725 (.Y (nx2724), .A0 (nx2662), .A1 (nx1805), .S0 (nx2666)) ;
    xnor2 ix2663 (.Y (nx2662), .A0 (nx1743), .A1 (nx2326)) ;
    mux21 ix1806 (.Y (nx1805), .A0 (nx1807), .A1 (nx2716), .S0 (nx2678)) ;
    xnor2 ix1808 (.Y (nx1807), .A0 (nx2356), .A1 (nx2334)) ;
    mux21 ix2717 (.Y (nx2716), .A0 (nx2686), .A1 (nx1813), .S0 (nx2690)) ;
    xnor2 ix2687 (.Y (nx2686), .A0 (nx1755), .A1 (nx2346)) ;
    nor02ii ix1814 (.Y (nx1813), .A0 (nx1815), .A1 (nx1817)) ;
    oai21 ix1816 (.Y (nx1815), .A0 (T02[0]), .A1 (T22[0]), .B0 (nx1755)) ;
    oai21 ix1818 (.Y (nx1817), .A0 (T20[0]), .A1 (T00[0]), .B0 (nx1819)) ;
    nand02 ix1820 (.Y (nx1819), .A0 (T00[0]), .A1 (T20[0])) ;
    xnor2 ix2691 (.Y (nx2690), .A0 (nx2688), .A1 (nx2686)) ;
    xnor2 ix2689 (.Y (nx2688), .A0 (nx1819), .A1 (nx2510)) ;
    xnor2 ix2511 (.Y (nx2510), .A0 (T20[1]), .A1 (nx1827)) ;
    oai21 ix1828 (.Y (nx1827), .A0 (T10[0]), .A1 (T00[1]), .B0 (nx1829)) ;
    nand02 ix1830 (.Y (nx1829), .A0 (T00[1]), .A1 (T10[0])) ;
    xnor2 ix2679 (.Y (nx2678), .A0 (nx1833), .A1 (nx1807)) ;
    xnor2 ix1834 (.Y (nx1833), .A0 (nx2520), .A1 (nx2498)) ;
    mux21 ix2521 (.Y (nx2520), .A0 (nx1827), .A1 (nx1819), .S0 (nx2510)) ;
    xnor2 ix2499 (.Y (nx2498), .A0 (T20[2]), .A1 (nx1839)) ;
    xnor2 ix1840 (.Y (nx1839), .A0 (nx1829), .A1 (nx1841)) ;
    xnor2 ix1842 (.Y (nx1841), .A0 (T00[2]), .A1 (T10[1])) ;
    xnor2 ix2667 (.Y (nx2666), .A0 (nx2664), .A1 (nx2662)) ;
    xnor2 ix2665 (.Y (nx2664), .A0 (nx1847), .A1 (nx2490)) ;
    aoi22 ix1848 (.Y (nx1847), .A0 (nx2496), .A1 (T20[2]), .B0 (nx2520), .B1 (
          nx2498)) ;
    xnor2 ix2491 (.Y (nx2490), .A0 (T20[3]), .A1 (nx1853)) ;
    xnor2 ix1854 (.Y (nx1853), .A0 (nx1855), .A1 (nx1861)) ;
    aoi32 ix1856 (.Y (nx1855), .A0 (T00[1]), .A1 (T10[0]), .A2 (nx2426), .B0 (
          T10[1]), .B1 (T00[2])) ;
    xnor2 ix1862 (.Y (nx1861), .A0 (T00[3]), .A1 (T10[2])) ;
    xnor2 ix2655 (.Y (nx2654), .A0 (nx2652), .A1 (nx2650)) ;
    xnor2 ix2653 (.Y (nx2652), .A0 (nx2528), .A1 (nx1869)) ;
    mux21 ix2529 (.Y (nx2528), .A0 (nx1853), .A1 (nx1847), .S0 (nx2490)) ;
    xnor2 ix1870 (.Y (nx1869), .A0 (T20[4]), .A1 (nx2480)) ;
    xnor2 ix2481 (.Y (nx2480), .A0 (nx2440), .A1 (nx1877)) ;
    mux21 ix2441 (.Y (nx2440), .A0 (nx1855), .A1 (nx1875), .S0 (nx1861)) ;
    inv01 ix1876 (.Y (nx1875), .A (T10[2])) ;
    xnor2 ix1878 (.Y (nx1877), .A0 (T00[4]), .A1 (T10[3])) ;
    xnor2 ix2651 (.Y (nx2650), .A0 (nx2364), .A1 (nx1767)) ;
    xnor2 ix2643 (.Y (nx2642), .A0 (nx2640), .A1 (nx2638)) ;
    xnor2 ix2641 (.Y (nx2640), .A0 (nx1885), .A1 (nx2474)) ;
    mux21 ix1886 (.Y (nx1885), .A0 (nx2528), .A1 (nx2480), .S0 (nx1869)) ;
    xnor2 ix2475 (.Y (nx2474), .A0 (T20[5]), .A1 (nx1889)) ;
    xnor2 ix1890 (.Y (nx1889), .A0 (nx1891), .A1 (nx1893)) ;
    mux21 ix1892 (.Y (nx1891), .A0 (nx2440), .A1 (T10[3]), .S0 (nx1877)) ;
    xnor2 ix1894 (.Y (nx1893), .A0 (T00[5]), .A1 (T10[4])) ;
    xnor2 ix2631 (.Y (nx2630), .A0 (nx2628), .A1 (nx2626)) ;
    xnor2 ix2629 (.Y (nx2628), .A0 (nx2536), .A1 (nx1901)) ;
    mux21 ix2537 (.Y (nx2536), .A0 (nx1889), .A1 (nx1885), .S0 (nx2474)) ;
    xnor2 ix1902 (.Y (nx1901), .A0 (T20[6]), .A1 (nx2464)) ;
    xnor2 ix2465 (.Y (nx2464), .A0 (nx2448), .A1 (nx1909)) ;
    mux21 ix2449 (.Y (nx2448), .A0 (nx1891), .A1 (nx1907), .S0 (nx1893)) ;
    inv01 ix1908 (.Y (nx1907), .A (T10[4])) ;
    xnor2 ix1910 (.Y (nx1909), .A0 (T00[6]), .A1 (T10[5])) ;
    xnor2 ix2627 (.Y (nx2626), .A0 (nx2372), .A1 (nx1773)) ;
    xnor2 ix2619 (.Y (nx2618), .A0 (nx2616), .A1 (nx2614)) ;
    xnor2 ix2617 (.Y (nx2616), .A0 (nx1917), .A1 (nx2458)) ;
    mux21 ix1918 (.Y (nx1917), .A0 (nx2536), .A1 (nx2464), .S0 (nx1901)) ;
    xnor2 ix2459 (.Y (nx2458), .A0 (T20[7]), .A1 (nx1921)) ;
    xnor2 ix1922 (.Y (nx1921), .A0 (nx1923), .A1 (nx1925)) ;
    mux21 ix1924 (.Y (nx1923), .A0 (nx2448), .A1 (T10[5]), .S0 (nx1909)) ;
    xnor2 ix1926 (.Y (nx1925), .A0 (T00[7]), .A1 (T10[6])) ;
    xnor2 ix2607 (.Y (nx2606), .A0 (nx2604), .A1 (nx2598)) ;
    xnor2 ix2605 (.Y (nx2604), .A0 (nx2544), .A1 (nx1933)) ;
    mux21 ix2545 (.Y (nx2544), .A0 (nx1921), .A1 (nx1917), .S0 (nx2458)) ;
    xnor2 ix1934 (.Y (nx1933), .A0 (T10[7]), .A1 (nx2552)) ;
    mux21 ix2553 (.Y (nx2552), .A0 (nx1923), .A1 (nx1937), .S0 (nx1925)) ;
    inv01 ix1938 (.Y (nx1937), .A (T10[6])) ;
    xnor2 ix2599 (.Y (nx2598), .A0 (nx2380), .A1 (nx1783)) ;
    xnor2 ix2587 (.Y (nx2586), .A0 (nx1943), .A1 (nx1951)) ;
    nor02ii ix1946 (.Y (nx1943), .A0 (nx2562), .A1 (nx1949)) ;
    nor02ii ix2563 (.Y (nx2562), .A0 (nx1933), .A1 (nx2544)) ;
    nand02 ix1950 (.Y (nx1949), .A0 (T10[7]), .A1 (nx2552)) ;
    nor02ii ix1954 (.Y (nx1951), .A0 (nx2398), .A1 (nx1691)) ;
    nor02ii ix2399 (.Y (nx2398), .A0 (nx1783), .A1 (nx2380)) ;
    mux21 ix1958 (.Y (nx1957), .A0 (nx2852), .A1 (nx3182), .S0 (nx2447)) ;
    mux21 ix2847 (.Y (nx2846), .A0 (nx2580), .A1 (nx1969), .S0 (nx2586)) ;
    mux21 ix1970 (.Y (nx1969), .A0 (nx1971), .A1 (nx2838), .S0 (nx2606)) ;
    mux21 ix2839 (.Y (nx2838), .A0 (nx2616), .A1 (nx1975), .S0 (nx2618)) ;
    mux21 ix1976 (.Y (nx1975), .A0 (nx1977), .A1 (nx2830), .S0 (nx2630)) ;
    mux21 ix2831 (.Y (nx2830), .A0 (nx2640), .A1 (nx1981), .S0 (nx2642)) ;
    mux21 ix1982 (.Y (nx1981), .A0 (nx1983), .A1 (nx2822), .S0 (nx2654)) ;
    mux21 ix2823 (.Y (nx2822), .A0 (nx2664), .A1 (nx1987), .S0 (nx2666)) ;
    mux21 ix1988 (.Y (nx1987), .A0 (nx1833), .A1 (nx2814), .S0 (nx2678)) ;
    mux21 ix2815 (.Y (nx2814), .A0 (nx2688), .A1 (nx1991), .S0 (nx2690)) ;
    nor02ii ix1992 (.Y (nx1991), .A0 (nx1817), .A1 (nx1815)) ;
    mux21 ix3183 (.Y (nx3182), .A0 (nx1995), .A1 (nx2007), .S0 (nx2435)) ;
    xnor2 ix2869 (.Y (nx2868), .A0 (nx1779), .A1 (nx2586)) ;
    xnor2 ix2863 (.Y (nx2862), .A0 (nx1969), .A1 (nx2586)) ;
    nand02 ix2004 (.Y (nx2001), .A0 (nx2748), .A1 (nx360)) ;
    mux21 ix2008 (.Y (nx2007), .A0 (nx2898), .A1 (nx3166), .S0 (nx2425)) ;
    xnor2 ix2012 (.Y (nx2011), .A0 (nx2740), .A1 (nx2606)) ;
    xnor2 ix2014 (.Y (nx2013), .A0 (nx2838), .A1 (nx2606)) ;
    mux21 ix3167 (.Y (nx3166), .A0 (nx2017), .A1 (nx2023), .S0 (nx2413)) ;
    xnor2 ix2921 (.Y (nx2920), .A0 (nx1789), .A1 (nx2618)) ;
    xnor2 ix2915 (.Y (nx2914), .A0 (nx1975), .A1 (nx2618)) ;
    mux21 ix2024 (.Y (nx2023), .A0 (nx2950), .A1 (nx3150), .S0 (nx2403)) ;
    xnor2 ix2028 (.Y (nx2027), .A0 (nx2732), .A1 (nx2630)) ;
    xnor2 ix2030 (.Y (nx2029), .A0 (nx2830), .A1 (nx2630)) ;
    mux21 ix3151 (.Y (nx3150), .A0 (nx2033), .A1 (nx2039), .S0 (nx2391)) ;
    xnor2 ix2973 (.Y (nx2972), .A0 (nx1797), .A1 (nx2642)) ;
    xnor2 ix2967 (.Y (nx2966), .A0 (nx1981), .A1 (nx2642)) ;
    mux21 ix2040 (.Y (nx2039), .A0 (nx3002), .A1 (nx3134), .S0 (nx2381)) ;
    xnor2 ix2044 (.Y (nx2043), .A0 (nx2724), .A1 (nx2654)) ;
    xnor2 ix2046 (.Y (nx2045), .A0 (nx2822), .A1 (nx2654)) ;
    mux21 ix3135 (.Y (nx3134), .A0 (nx2049), .A1 (nx2055), .S0 (nx2371)) ;
    xnor2 ix3025 (.Y (nx3024), .A0 (nx1805), .A1 (nx2666)) ;
    xnor2 ix3019 (.Y (nx3018), .A0 (nx1987), .A1 (nx2666)) ;
    mux21 ix2056 (.Y (nx2055), .A0 (nx3054), .A1 (nx3118), .S0 (nx2361)) ;
    xnor2 ix2060 (.Y (nx2059), .A0 (nx2716), .A1 (nx2678)) ;
    xnor2 ix2062 (.Y (nx2061), .A0 (nx2814), .A1 (nx2678)) ;
    mux21 ix3119 (.Y (nx3118), .A0 (nx2065), .A1 (nx2071), .S0 (nx2089)) ;
    xnor2 ix3077 (.Y (nx3076), .A0 (nx1813), .A1 (nx2690)) ;
    xnor2 ix3071 (.Y (nx3070), .A0 (nx1991), .A1 (nx2690)) ;
    nand02 ix2072 (.Y (nx2071), .A0 (nx3100), .A1 (nx2075)) ;
    nor02 ix2076 (.Y (nx2075), .A0 (nx2077), .A1 (nx2087)) ;
    nor02ii ix2078 (.Y (nx2077), .A0 (nx2079), .A1 (nx2083)) ;
    oai21 ix2080 (.Y (nx2079), .A0 (T12[0]), .A1 (T21[0]), .B0 (nx2081)) ;
    nand02 ix2082 (.Y (nx2081), .A0 (T21[0]), .A1 (T12[0])) ;
    oai21 ix2084 (.Y (nx2083), .A0 (T01[0]), .A1 (T10[0]), .B0 (nx2085)) ;
    nand02 ix2086 (.Y (nx2085), .A0 (T10[0]), .A1 (T01[0])) ;
    nor02ii ix2088 (.Y (nx2087), .A0 (nx2083), .A1 (nx2079)) ;
    xnor2 ix2090 (.Y (nx2089), .A0 (nx2065), .A1 (nx2091)) ;
    xnor2 ix3089 (.Y (nx3088), .A0 (nx2087), .A1 (nx2068)) ;
    xnor2 ix2069 (.Y (nx2068), .A0 (nx2066), .A1 (nx2064)) ;
    xnor2 ix2067 (.Y (nx2066), .A0 (nx2081), .A1 (nx1888)) ;
    xnor2 ix1889 (.Y (nx1888), .A0 (T12[1]), .A1 (nx2101)) ;
    oai21 ix2102 (.Y (nx2101), .A0 (T21[1]), .A1 (T22[0]), .B0 (nx2103)) ;
    nand02 ix2104 (.Y (nx2103), .A0 (T22[0]), .A1 (T21[1])) ;
    xnor2 ix2065 (.Y (nx2064), .A0 (nx2085), .A1 (nx1724)) ;
    xnor2 ix1725 (.Y (nx1724), .A0 (T01[1]), .A1 (nx2109)) ;
    oai21 ix2110 (.Y (nx2109), .A0 (T10[1]), .A1 (T00[0]), .B0 (nx2111)) ;
    nand02 ix2112 (.Y (nx2111), .A0 (T00[0]), .A1 (T10[1])) ;
    xnor2 ix3083 (.Y (nx3082), .A0 (nx2077), .A1 (nx2068)) ;
    nand02 ix2118 (.Y (nx2115), .A0 (nx2126), .A1 (nx360)) ;
    mux21 ix2127 (.Y (nx2126), .A0 (nx1952), .A1 (nx2201), .S0 (nx1964)) ;
    nand02 ix2124 (.Y (nx2123), .A0 (T00[7]), .A1 (nx1766)) ;
    mux21 ix1767 (.Y (nx1766), .A0 (nx2127), .A1 (nx2151), .S0 (nx2153)) ;
    mux21 ix2128 (.Y (nx2127), .A0 (nx1662), .A1 (T10[6]), .S0 (nx2149)) ;
    mux21 ix1663 (.Y (nx1662), .A0 (nx2131), .A1 (nx2145), .S0 (nx2147)) ;
    mux21 ix2132 (.Y (nx2131), .A0 (nx1654), .A1 (T10[4]), .S0 (nx2143)) ;
    mux21 ix1655 (.Y (nx1654), .A0 (nx2135), .A1 (nx2139), .S0 (nx2141)) ;
    aoi32 ix2136 (.Y (nx2135), .A0 (T00[0]), .A1 (T10[1]), .A2 (nx1640), .B0 (
          T10[2]), .B1 (T00[1])) ;
    inv01 ix2140 (.Y (nx2139), .A (T10[3])) ;
    xnor2 ix2142 (.Y (nx2141), .A0 (T00[2]), .A1 (T10[3])) ;
    xnor2 ix2144 (.Y (nx2143), .A0 (T00[3]), .A1 (T10[4])) ;
    inv01 ix2146 (.Y (nx2145), .A (T10[5])) ;
    xnor2 ix2148 (.Y (nx2147), .A0 (T00[4]), .A1 (T10[5])) ;
    xnor2 ix2150 (.Y (nx2149), .A0 (T00[5]), .A1 (T10[6])) ;
    inv01 ix2152 (.Y (nx2151), .A (T10[7])) ;
    xnor2 ix2154 (.Y (nx2153), .A0 (T00[6]), .A1 (T10[7])) ;
    mux21 ix1759 (.Y (nx1758), .A0 (nx2159), .A1 (nx2161), .S0 (nx1672)) ;
    xnor2 ix2160 (.Y (nx2159), .A0 (nx2127), .A1 (nx2153)) ;
    mux21 ix2162 (.Y (nx2161), .A0 (nx1750), .A1 (nx1678), .S0 (nx2195)) ;
    mux21 ix1751 (.Y (nx1750), .A0 (nx2165), .A1 (nx2167), .S0 (nx1688)) ;
    xnor2 ix2166 (.Y (nx2165), .A0 (nx2131), .A1 (nx2147)) ;
    mux21 ix2168 (.Y (nx2167), .A0 (nx1742), .A1 (nx1694), .S0 (nx2189)) ;
    mux21 ix1743 (.Y (nx1742), .A0 (nx2171), .A1 (nx2173), .S0 (nx1704)) ;
    xnor2 ix2172 (.Y (nx2171), .A0 (nx2135), .A1 (nx2141)) ;
    aoi22 ix2174 (.Y (nx2173), .A0 (nx1710), .A1 (T01[2]), .B0 (nx1734), .B1 (
          nx1712)) ;
    xnor2 ix2178 (.Y (nx2177), .A0 (T00[1]), .A1 (T10[2])) ;
    mux21 ix1735 (.Y (nx1734), .A0 (nx2109), .A1 (nx2085), .S0 (nx1724)) ;
    xnor2 ix1713 (.Y (nx1712), .A0 (T01[2]), .A1 (nx2183)) ;
    xnor2 ix2184 (.Y (nx2183), .A0 (nx2111), .A1 (nx2177)) ;
    xnor2 ix1705 (.Y (nx1704), .A0 (T01[3]), .A1 (nx2171)) ;
    xnor2 ix1695 (.Y (nx1694), .A0 (nx1654), .A1 (nx2143)) ;
    xnor2 ix2190 (.Y (nx2189), .A0 (T01[4]), .A1 (nx1694)) ;
    xnor2 ix1689 (.Y (nx1688), .A0 (T01[5]), .A1 (nx2165)) ;
    xnor2 ix1679 (.Y (nx1678), .A0 (nx1662), .A1 (nx2149)) ;
    xnor2 ix2196 (.Y (nx2195), .A0 (T01[6]), .A1 (nx1678)) ;
    xnor2 ix1673 (.Y (nx1672), .A0 (T01[7]), .A1 (nx2159)) ;
    mux21 ix2202 (.Y (nx2201), .A0 (nx2203), .A1 (nx2118), .S0 (nx1984)) ;
    xnor2 ix2206 (.Y (nx2205), .A0 (T00[7]), .A1 (nx1766)) ;
    mux21 ix2119 (.Y (nx2118), .A0 (nx1992), .A1 (nx2211), .S0 (nx1996)) ;
    xnor2 ix1993 (.Y (nx1992), .A0 (nx2161), .A1 (nx1672)) ;
    mux21 ix2212 (.Y (nx2211), .A0 (nx2213), .A1 (nx2110), .S0 (nx2008)) ;
    mux21 ix2111 (.Y (nx2110), .A0 (nx2016), .A1 (nx2219), .S0 (nx2020)) ;
    xnor2 ix2017 (.Y (nx2016), .A0 (nx2167), .A1 (nx1688)) ;
    mux21 ix2220 (.Y (nx2219), .A0 (nx2221), .A1 (nx2102), .S0 (nx2032)) ;
    mux21 ix2103 (.Y (nx2102), .A0 (nx2040), .A1 (nx2227), .S0 (nx2044)) ;
    xnor2 ix2041 (.Y (nx2040), .A0 (nx2173), .A1 (nx1704)) ;
    mux21 ix2228 (.Y (nx2227), .A0 (nx2229), .A1 (nx2094), .S0 (nx2056)) ;
    xnor2 ix2230 (.Y (nx2229), .A0 (nx1734), .A1 (nx1712)) ;
    mux21 ix2095 (.Y (nx2094), .A0 (nx2064), .A1 (nx2087), .S0 (nx2068)) ;
    xnor2 ix2057 (.Y (nx2056), .A0 (nx2235), .A1 (nx2229)) ;
    xnor2 ix2236 (.Y (nx2235), .A0 (nx1898), .A1 (nx1876)) ;
    mux21 ix1899 (.Y (nx1898), .A0 (nx2101), .A1 (nx2081), .S0 (nx1888)) ;
    xnor2 ix1877 (.Y (nx1876), .A0 (T12[2]), .A1 (nx2241)) ;
    xnor2 ix2242 (.Y (nx2241), .A0 (nx2103), .A1 (nx2243)) ;
    xnor2 ix2244 (.Y (nx2243), .A0 (T22[1]), .A1 (T21[2])) ;
    xnor2 ix2045 (.Y (nx2044), .A0 (nx2042), .A1 (nx2040)) ;
    xnor2 ix2043 (.Y (nx2042), .A0 (nx2249), .A1 (nx1868)) ;
    aoi22 ix2250 (.Y (nx2249), .A0 (nx1874), .A1 (T12[2]), .B0 (nx1898), .B1 (
          nx1876)) ;
    xnor2 ix1869 (.Y (nx1868), .A0 (T12[3]), .A1 (nx2255)) ;
    xnor2 ix2256 (.Y (nx2255), .A0 (nx2257), .A1 (nx2263)) ;
    aoi32 ix2258 (.Y (nx2257), .A0 (T22[0]), .A1 (T21[1]), .A2 (nx1804), .B0 (
          T21[2]), .B1 (T22[1])) ;
    xnor2 ix2264 (.Y (nx2263), .A0 (T22[2]), .A1 (T21[3])) ;
    xnor2 ix2033 (.Y (nx2032), .A0 (nx2030), .A1 (nx2028)) ;
    xnor2 ix2031 (.Y (nx2030), .A0 (nx1906), .A1 (nx2271)) ;
    mux21 ix1907 (.Y (nx1906), .A0 (nx2255), .A1 (nx2249), .S0 (nx1868)) ;
    xnor2 ix2272 (.Y (nx2271), .A0 (T12[4]), .A1 (nx1858)) ;
    xnor2 ix1859 (.Y (nx1858), .A0 (nx1818), .A1 (nx2279)) ;
    mux21 ix1819 (.Y (nx1818), .A0 (nx2257), .A1 (nx2277), .S0 (nx2263)) ;
    inv01 ix2278 (.Y (nx2277), .A (T21[3])) ;
    xnor2 ix2280 (.Y (nx2279), .A0 (T22[3]), .A1 (T21[4])) ;
    xnor2 ix2029 (.Y (nx2028), .A0 (nx1742), .A1 (nx2189)) ;
    xnor2 ix2021 (.Y (nx2020), .A0 (nx2018), .A1 (nx2016)) ;
    xnor2 ix2019 (.Y (nx2018), .A0 (nx2287), .A1 (nx1852)) ;
    mux21 ix2288 (.Y (nx2287), .A0 (nx1906), .A1 (nx1858), .S0 (nx2271)) ;
    xnor2 ix1853 (.Y (nx1852), .A0 (T12[5]), .A1 (nx2291)) ;
    xnor2 ix2292 (.Y (nx2291), .A0 (nx2293), .A1 (nx2295)) ;
    mux21 ix2294 (.Y (nx2293), .A0 (nx1818), .A1 (T21[4]), .S0 (nx2279)) ;
    xnor2 ix2296 (.Y (nx2295), .A0 (T22[4]), .A1 (T21[5])) ;
    xnor2 ix2009 (.Y (nx2008), .A0 (nx2006), .A1 (nx2004)) ;
    xnor2 ix2007 (.Y (nx2006), .A0 (nx1914), .A1 (nx2303)) ;
    mux21 ix1915 (.Y (nx1914), .A0 (nx2291), .A1 (nx2287), .S0 (nx1852)) ;
    xnor2 ix2304 (.Y (nx2303), .A0 (T12[6]), .A1 (nx1842)) ;
    xnor2 ix1843 (.Y (nx1842), .A0 (nx1826), .A1 (nx2311)) ;
    mux21 ix1827 (.Y (nx1826), .A0 (nx2293), .A1 (nx2309), .S0 (nx2295)) ;
    inv01 ix2310 (.Y (nx2309), .A (T21[5])) ;
    xnor2 ix2312 (.Y (nx2311), .A0 (T22[5]), .A1 (T21[6])) ;
    xnor2 ix2005 (.Y (nx2004), .A0 (nx1750), .A1 (nx2195)) ;
    xnor2 ix1997 (.Y (nx1996), .A0 (nx1994), .A1 (nx1992)) ;
    xnor2 ix1995 (.Y (nx1994), .A0 (nx2319), .A1 (nx1836)) ;
    mux21 ix2320 (.Y (nx2319), .A0 (nx1914), .A1 (nx1842), .S0 (nx2303)) ;
    xnor2 ix1837 (.Y (nx1836), .A0 (T12[7]), .A1 (nx2323)) ;
    xnor2 ix2324 (.Y (nx2323), .A0 (nx2325), .A1 (nx2327)) ;
    mux21 ix2326 (.Y (nx2325), .A0 (nx1826), .A1 (T21[6]), .S0 (nx2311)) ;
    xnor2 ix2328 (.Y (nx2327), .A0 (T22[6]), .A1 (T21[7])) ;
    xnor2 ix1985 (.Y (nx1984), .A0 (nx1982), .A1 (nx1976)) ;
    xnor2 ix1983 (.Y (nx1982), .A0 (nx1922), .A1 (nx2335)) ;
    mux21 ix1923 (.Y (nx1922), .A0 (nx2323), .A1 (nx2319), .S0 (nx1836)) ;
    xnor2 ix2336 (.Y (nx2335), .A0 (T22[7]), .A1 (nx1930)) ;
    mux21 ix1931 (.Y (nx1930), .A0 (nx2325), .A1 (nx2339), .S0 (nx2327)) ;
    inv01 ix2340 (.Y (nx2339), .A (T21[7])) ;
    xnor2 ix1977 (.Y (nx1976), .A0 (nx1758), .A1 (nx2205)) ;
    xnor2 ix1965 (.Y (nx1964), .A0 (nx2345), .A1 (nx2353)) ;
    nor02ii ix2348 (.Y (nx2345), .A0 (nx1940), .A1 (nx2351)) ;
    nor02ii ix1941 (.Y (nx1940), .A0 (nx2335), .A1 (nx1922)) ;
    nand02 ix2352 (.Y (nx2351), .A0 (T22[7]), .A1 (nx1930)) ;
    nor02ii ix2356 (.Y (nx2353), .A0 (nx1776), .A1 (nx2123)) ;
    nor02ii ix1777 (.Y (nx1776), .A0 (nx2205), .A1 (nx1758)) ;
    xnor2 ix2362 (.Y (nx2361), .A0 (nx3054), .A1 (nx3066)) ;
    xnor2 ix2366 (.Y (nx2365), .A0 (nx2094), .A1 (nx2056)) ;
    xnor2 ix2368 (.Y (nx2367), .A0 (nx2192), .A1 (nx2056)) ;
    mux21 ix2193 (.Y (nx2192), .A0 (nx2066), .A1 (nx2077), .S0 (nx2068)) ;
    xnor2 ix2372 (.Y (nx2371), .A0 (nx2049), .A1 (nx2373)) ;
    xnor2 ix3037 (.Y (nx3036), .A0 (nx2227), .A1 (nx2044)) ;
    xnor2 ix3031 (.Y (nx3030), .A0 (nx2379), .A1 (nx2044)) ;
    mux21 ix2380 (.Y (nx2379), .A0 (nx2235), .A1 (nx2192), .S0 (nx2056)) ;
    xnor2 ix2382 (.Y (nx2381), .A0 (nx3002), .A1 (nx3014)) ;
    xnor2 ix2386 (.Y (nx2385), .A0 (nx2102), .A1 (nx2032)) ;
    xnor2 ix2388 (.Y (nx2387), .A0 (nx2200), .A1 (nx2032)) ;
    mux21 ix2201 (.Y (nx2200), .A0 (nx2042), .A1 (nx2379), .S0 (nx2044)) ;
    xnor2 ix2392 (.Y (nx2391), .A0 (nx2033), .A1 (nx2393)) ;
    xnor2 ix2985 (.Y (nx2984), .A0 (nx2219), .A1 (nx2020)) ;
    xnor2 ix2979 (.Y (nx2978), .A0 (nx2399), .A1 (nx2020)) ;
    mux21 ix2400 (.Y (nx2399), .A0 (nx2401), .A1 (nx2200), .S0 (nx2032)) ;
    xnor2 ix2404 (.Y (nx2403), .A0 (nx2950), .A1 (nx2962)) ;
    xnor2 ix2408 (.Y (nx2407), .A0 (nx2110), .A1 (nx2008)) ;
    xnor2 ix2410 (.Y (nx2409), .A0 (nx2208), .A1 (nx2008)) ;
    mux21 ix2209 (.Y (nx2208), .A0 (nx2018), .A1 (nx2399), .S0 (nx2020)) ;
    xnor2 ix2414 (.Y (nx2413), .A0 (nx2017), .A1 (nx2415)) ;
    xnor2 ix2933 (.Y (nx2932), .A0 (nx2211), .A1 (nx1996)) ;
    xnor2 ix2927 (.Y (nx2926), .A0 (nx2421), .A1 (nx1996)) ;
    mux21 ix2422 (.Y (nx2421), .A0 (nx2423), .A1 (nx2208), .S0 (nx2008)) ;
    xnor2 ix2426 (.Y (nx2425), .A0 (nx2898), .A1 (nx2910)) ;
    xnor2 ix2430 (.Y (nx2429), .A0 (nx2118), .A1 (nx1984)) ;
    xnor2 ix2432 (.Y (nx2431), .A0 (nx2216), .A1 (nx1984)) ;
    mux21 ix2217 (.Y (nx2216), .A0 (nx1994), .A1 (nx2421), .S0 (nx1996)) ;
    xnor2 ix2436 (.Y (nx2435), .A0 (nx1995), .A1 (nx2437)) ;
    xnor2 ix2881 (.Y (nx2880), .A0 (nx2201), .A1 (nx1964)) ;
    xnor2 ix2875 (.Y (nx2874), .A0 (nx2443), .A1 (nx1964)) ;
    mux21 ix2444 (.Y (nx2443), .A0 (nx2445), .A1 (nx2216), .S0 (nx1984)) ;
    xnor2 ix2448 (.Y (nx2447), .A0 (nx2852), .A1 (nx2230)) ;
    mux21 ix2225 (.Y (nx2224), .A0 (nx1958), .A1 (nx2443), .S0 (nx1964)) ;
    mux21 ix3463 (.Y (nx3462), .A0 (nx2465), .A1 (nx3055), .S0 (nx3299)) ;
    nor02 ix2466 (.Y (nx2465), .A0 (nx646), .A1 (nx1268)) ;
    mux21 ix543 (.Y (nx542), .A0 (nx368), .A1 (nx2563), .S0 (nx380)) ;
    nand02 ix2476 (.Y (nx2475), .A0 (T02[7]), .A1 (nx182)) ;
    mux21 ix183 (.Y (nx182), .A0 (nx2479), .A1 (nx2505), .S0 (nx2507)) ;
    mux21 ix2480 (.Y (nx2479), .A0 (nx78), .A1 (T01[6]), .S0 (nx2503)) ;
    mux21 ix79 (.Y (nx78), .A0 (nx2483), .A1 (nx2499), .S0 (nx2501)) ;
    mux21 ix2484 (.Y (nx2483), .A0 (nx70), .A1 (T01[4]), .S0 (nx2497)) ;
    mux21 ix71 (.Y (nx70), .A0 (nx2487), .A1 (nx2493), .S0 (nx2495)) ;
    aoi32 ix2488 (.Y (nx2487), .A0 (T02[0]), .A1 (T01[1]), .A2 (nx56), .B0 (
          T01[2]), .B1 (T02[1])) ;
    inv01 ix2492 (.Y (nx2491), .A (T01[2])) ;
    inv01 ix2494 (.Y (nx2493), .A (T01[3])) ;
    xnor2 ix2496 (.Y (nx2495), .A0 (T02[2]), .A1 (T01[3])) ;
    xnor2 ix2498 (.Y (nx2497), .A0 (T02[3]), .A1 (T01[4])) ;
    inv01 ix2500 (.Y (nx2499), .A (T01[5])) ;
    xnor2 ix2502 (.Y (nx2501), .A0 (T02[4]), .A1 (T01[5])) ;
    xnor2 ix2504 (.Y (nx2503), .A0 (T02[5]), .A1 (T01[6])) ;
    inv01 ix2506 (.Y (nx2505), .A (T01[7])) ;
    xnor2 ix2508 (.Y (nx2507), .A0 (T02[6]), .A1 (T01[7])) ;
    mux21 ix175 (.Y (nx174), .A0 (nx2513), .A1 (nx2515), .S0 (nx88)) ;
    xnor2 ix2514 (.Y (nx2513), .A0 (nx2479), .A1 (nx2507)) ;
    mux21 ix2516 (.Y (nx2515), .A0 (nx166), .A1 (nx94), .S0 (nx2557)) ;
    mux21 ix167 (.Y (nx166), .A0 (nx2519), .A1 (nx2521), .S0 (nx104)) ;
    xnor2 ix2520 (.Y (nx2519), .A0 (nx2483), .A1 (nx2501)) ;
    mux21 ix2522 (.Y (nx2521), .A0 (nx158), .A1 (nx110), .S0 (nx2551)) ;
    mux21 ix159 (.Y (nx158), .A0 (nx2525), .A1 (nx2527), .S0 (nx120)) ;
    xnor2 ix2526 (.Y (nx2525), .A0 (nx2487), .A1 (nx2495)) ;
    aoi22 ix2528 (.Y (nx2527), .A0 (nx126), .A1 (T12[2]), .B0 (nx150), .B1 (
          nx128)) ;
    nand02 ix2532 (.Y (nx2531), .A0 (T02[0]), .A1 (T01[1])) ;
    xnor2 ix2534 (.Y (nx2533), .A0 (T02[1]), .A1 (T01[2])) ;
    mux21 ix151 (.Y (nx150), .A0 (nx2537), .A1 (nx2539), .S0 (nx140)) ;
    oai21 ix2538 (.Y (nx2537), .A0 (T01[1]), .A1 (T02[0]), .B0 (nx2531)) ;
    nand02 ix2540 (.Y (nx2539), .A0 (T12[0]), .A1 (T01[0])) ;
    xnor2 ix141 (.Y (nx140), .A0 (T12[1]), .A1 (nx2537)) ;
    xnor2 ix129 (.Y (nx128), .A0 (T12[2]), .A1 (nx2545)) ;
    xnor2 ix2546 (.Y (nx2545), .A0 (nx2531), .A1 (nx2533)) ;
    xnor2 ix121 (.Y (nx120), .A0 (T12[3]), .A1 (nx2525)) ;
    xnor2 ix111 (.Y (nx110), .A0 (nx70), .A1 (nx2497)) ;
    xnor2 ix2552 (.Y (nx2551), .A0 (T12[4]), .A1 (nx110)) ;
    xnor2 ix105 (.Y (nx104), .A0 (T12[5]), .A1 (nx2519)) ;
    xnor2 ix95 (.Y (nx94), .A0 (nx78), .A1 (nx2503)) ;
    xnor2 ix2558 (.Y (nx2557), .A0 (T12[6]), .A1 (nx94)) ;
    xnor2 ix89 (.Y (nx88), .A0 (T12[7]), .A1 (nx2513)) ;
    mux21 ix2564 (.Y (nx2563), .A0 (nx2565), .A1 (nx534), .S0 (nx400)) ;
    xnor2 ix2568 (.Y (nx2567), .A0 (T02[7]), .A1 (nx182)) ;
    mux21 ix535 (.Y (nx534), .A0 (nx408), .A1 (nx2573), .S0 (nx412)) ;
    xnor2 ix409 (.Y (nx408), .A0 (nx2515), .A1 (nx88)) ;
    mux21 ix2574 (.Y (nx2573), .A0 (nx2575), .A1 (nx526), .S0 (nx424)) ;
    mux21 ix527 (.Y (nx526), .A0 (nx432), .A1 (nx2579), .S0 (nx436)) ;
    xnor2 ix433 (.Y (nx432), .A0 (nx2521), .A1 (nx104)) ;
    mux21 ix2580 (.Y (nx2579), .A0 (nx2581), .A1 (nx518), .S0 (nx448)) ;
    mux21 ix519 (.Y (nx518), .A0 (nx456), .A1 (nx2587), .S0 (nx460)) ;
    xnor2 ix457 (.Y (nx456), .A0 (nx2527), .A1 (nx120)) ;
    mux21 ix2588 (.Y (nx2587), .A0 (nx2589), .A1 (nx510), .S0 (nx472)) ;
    xnor2 ix2590 (.Y (nx2589), .A0 (nx150), .A1 (nx128)) ;
    mux21 ix511 (.Y (nx510), .A0 (nx480), .A1 (nx2595), .S0 (nx484)) ;
    xnor2 ix481 (.Y (nx480), .A0 (nx2539), .A1 (nx140)) ;
    nor02ii ix2596 (.Y (nx2595), .A0 (nx2597), .A1 (nx2599)) ;
    oai21 ix2598 (.Y (nx2597), .A0 (T01[0]), .A1 (T12[0]), .B0 (nx2539)) ;
    oai21 ix2600 (.Y (nx2599), .A0 (T10[0]), .A1 (T21[0]), .B0 (nx2601)) ;
    nand02 ix2602 (.Y (nx2601), .A0 (T21[0]), .A1 (T10[0])) ;
    xnor2 ix485 (.Y (nx484), .A0 (nx482), .A1 (nx480)) ;
    xnor2 ix483 (.Y (nx482), .A0 (nx2601), .A1 (nx304)) ;
    xnor2 ix305 (.Y (nx304), .A0 (T21[1]), .A1 (nx2609)) ;
    oai21 ix2610 (.Y (nx2609), .A0 (T10[1]), .A1 (T20[0]), .B0 (nx2611)) ;
    nand02 ix2612 (.Y (nx2611), .A0 (T20[0]), .A1 (T10[1])) ;
    xnor2 ix473 (.Y (nx472), .A0 (nx2615), .A1 (nx2589)) ;
    xnor2 ix2616 (.Y (nx2615), .A0 (nx314), .A1 (nx292)) ;
    mux21 ix315 (.Y (nx314), .A0 (nx2609), .A1 (nx2601), .S0 (nx304)) ;
    xnor2 ix293 (.Y (nx292), .A0 (T21[2]), .A1 (nx2621)) ;
    xnor2 ix2622 (.Y (nx2621), .A0 (nx2611), .A1 (nx2623)) ;
    xnor2 ix2624 (.Y (nx2623), .A0 (T20[1]), .A1 (T10[2])) ;
    xnor2 ix461 (.Y (nx460), .A0 (nx458), .A1 (nx456)) ;
    xnor2 ix459 (.Y (nx458), .A0 (nx2629), .A1 (nx284)) ;
    aoi22 ix2630 (.Y (nx2629), .A0 (nx290), .A1 (T21[2]), .B0 (nx314), .B1 (
          nx292)) ;
    xnor2 ix285 (.Y (nx284), .A0 (T21[3]), .A1 (nx2635)) ;
    xnor2 ix2636 (.Y (nx2635), .A0 (nx2637), .A1 (nx2641)) ;
    aoi32 ix2638 (.Y (nx2637), .A0 (T20[0]), .A1 (T10[1]), .A2 (nx220), .B0 (
          T10[2]), .B1 (T20[1])) ;
    xnor2 ix2642 (.Y (nx2641), .A0 (T20[2]), .A1 (T10[3])) ;
    xnor2 ix449 (.Y (nx448), .A0 (nx446), .A1 (nx444)) ;
    xnor2 ix447 (.Y (nx446), .A0 (nx322), .A1 (nx2649)) ;
    mux21 ix323 (.Y (nx322), .A0 (nx2635), .A1 (nx2629), .S0 (nx284)) ;
    xnor2 ix2650 (.Y (nx2649), .A0 (T21[4]), .A1 (nx274)) ;
    xnor2 ix275 (.Y (nx274), .A0 (nx234), .A1 (nx2655)) ;
    mux21 ix235 (.Y (nx234), .A0 (nx2637), .A1 (nx2139), .S0 (nx2641)) ;
    xnor2 ix2656 (.Y (nx2655), .A0 (T20[3]), .A1 (T10[4])) ;
    xnor2 ix445 (.Y (nx444), .A0 (nx158), .A1 (nx2551)) ;
    xnor2 ix437 (.Y (nx436), .A0 (nx434), .A1 (nx432)) ;
    xnor2 ix435 (.Y (nx434), .A0 (nx2663), .A1 (nx268)) ;
    mux21 ix2664 (.Y (nx2663), .A0 (nx322), .A1 (nx274), .S0 (nx2649)) ;
    xnor2 ix269 (.Y (nx268), .A0 (T21[5]), .A1 (nx2667)) ;
    xnor2 ix2668 (.Y (nx2667), .A0 (nx2669), .A1 (nx2671)) ;
    mux21 ix2670 (.Y (nx2669), .A0 (nx234), .A1 (T10[4]), .S0 (nx2655)) ;
    xnor2 ix2672 (.Y (nx2671), .A0 (T20[4]), .A1 (T10[5])) ;
    xnor2 ix425 (.Y (nx424), .A0 (nx422), .A1 (nx420)) ;
    xnor2 ix423 (.Y (nx422), .A0 (nx330), .A1 (nx2679)) ;
    mux21 ix331 (.Y (nx330), .A0 (nx2667), .A1 (nx2663), .S0 (nx268)) ;
    xnor2 ix2680 (.Y (nx2679), .A0 (T21[6]), .A1 (nx258)) ;
    xnor2 ix259 (.Y (nx258), .A0 (nx242), .A1 (nx2685)) ;
    mux21 ix243 (.Y (nx242), .A0 (nx2669), .A1 (nx2145), .S0 (nx2671)) ;
    xnor2 ix2686 (.Y (nx2685), .A0 (T20[5]), .A1 (T10[6])) ;
    xnor2 ix421 (.Y (nx420), .A0 (nx166), .A1 (nx2557)) ;
    xnor2 ix413 (.Y (nx412), .A0 (nx410), .A1 (nx408)) ;
    xnor2 ix411 (.Y (nx410), .A0 (nx2693), .A1 (nx252)) ;
    mux21 ix2694 (.Y (nx2693), .A0 (nx330), .A1 (nx258), .S0 (nx2679)) ;
    xnor2 ix253 (.Y (nx252), .A0 (T21[7]), .A1 (nx2697)) ;
    xnor2 ix2698 (.Y (nx2697), .A0 (nx2699), .A1 (nx2701)) ;
    mux21 ix2700 (.Y (nx2699), .A0 (nx242), .A1 (T10[6]), .S0 (nx2685)) ;
    xnor2 ix2702 (.Y (nx2701), .A0 (T20[6]), .A1 (T10[7])) ;
    xnor2 ix401 (.Y (nx400), .A0 (nx398), .A1 (nx392)) ;
    xnor2 ix399 (.Y (nx398), .A0 (nx338), .A1 (nx2709)) ;
    mux21 ix339 (.Y (nx338), .A0 (nx2697), .A1 (nx2693), .S0 (nx252)) ;
    xnor2 ix2710 (.Y (nx2709), .A0 (T20[7]), .A1 (nx346)) ;
    mux21 ix347 (.Y (nx346), .A0 (nx2699), .A1 (nx2151), .S0 (nx2701)) ;
    xnor2 ix393 (.Y (nx392), .A0 (nx174), .A1 (nx2567)) ;
    xnor2 ix381 (.Y (nx380), .A0 (nx2717), .A1 (nx2725)) ;
    nor02ii ix2720 (.Y (nx2717), .A0 (nx356), .A1 (nx2723)) ;
    nor02ii ix357 (.Y (nx356), .A0 (nx2709), .A1 (nx338)) ;
    nand02 ix2724 (.Y (nx2723), .A0 (T20[7]), .A1 (nx346)) ;
    nor02ii ix2728 (.Y (nx2725), .A0 (nx192), .A1 (nx2475)) ;
    nor02ii ix193 (.Y (nx192), .A0 (nx2567), .A1 (nx174)) ;
    mux21 ix641 (.Y (nx640), .A0 (nx374), .A1 (nx2739), .S0 (nx380)) ;
    mux21 ix2740 (.Y (nx2739), .A0 (nx2741), .A1 (nx632), .S0 (nx400)) ;
    mux21 ix633 (.Y (nx632), .A0 (nx410), .A1 (nx2745), .S0 (nx412)) ;
    mux21 ix2746 (.Y (nx2745), .A0 (nx2747), .A1 (nx624), .S0 (nx424)) ;
    mux21 ix625 (.Y (nx624), .A0 (nx434), .A1 (nx2751), .S0 (nx436)) ;
    mux21 ix2752 (.Y (nx2751), .A0 (nx2753), .A1 (nx616), .S0 (nx448)) ;
    mux21 ix617 (.Y (nx616), .A0 (nx458), .A1 (nx2757), .S0 (nx460)) ;
    mux21 ix2758 (.Y (nx2757), .A0 (nx2615), .A1 (nx608), .S0 (nx472)) ;
    mux21 ix609 (.Y (nx608), .A0 (nx482), .A1 (nx2761), .S0 (nx484)) ;
    nor02ii ix2762 (.Y (nx2761), .A0 (nx2599), .A1 (nx2597)) ;
    mux21 ix1165 (.Y (nx1164), .A0 (nx990), .A1 (nx2855), .S0 (nx1002)) ;
    nand02 ix2770 (.Y (nx2769), .A0 (T01[7]), .A1 (nx804)) ;
    mux21 ix805 (.Y (nx804), .A0 (nx2773), .A1 (nx2797), .S0 (nx2799)) ;
    mux21 ix2774 (.Y (nx2773), .A0 (nx700), .A1 (T01[5]), .S0 (nx2795)) ;
    mux21 ix701 (.Y (nx700), .A0 (nx2777), .A1 (nx2791), .S0 (nx2793)) ;
    mux21 ix2778 (.Y (nx2777), .A0 (nx692), .A1 (T01[3]), .S0 (nx2789)) ;
    mux21 ix693 (.Y (nx692), .A0 (nx2781), .A1 (nx2491), .S0 (nx2787)) ;
    aoi32 ix2782 (.Y (nx2781), .A0 (T00[1]), .A1 (T01[0]), .A2 (nx678), .B0 (
          T01[1]), .B1 (T00[2])) ;
    xnor2 ix2788 (.Y (nx2787), .A0 (T00[3]), .A1 (T01[2])) ;
    xnor2 ix2790 (.Y (nx2789), .A0 (T00[4]), .A1 (T01[3])) ;
    inv01 ix2792 (.Y (nx2791), .A (T01[4])) ;
    xnor2 ix2794 (.Y (nx2793), .A0 (T00[5]), .A1 (T01[4])) ;
    xnor2 ix2796 (.Y (nx2795), .A0 (T00[6]), .A1 (T01[5])) ;
    inv01 ix2798 (.Y (nx2797), .A (T01[6])) ;
    xnor2 ix2800 (.Y (nx2799), .A0 (T00[7]), .A1 (T01[6])) ;
    mux21 ix797 (.Y (nx796), .A0 (nx2805), .A1 (nx2807), .S0 (nx710)) ;
    xnor2 ix2806 (.Y (nx2805), .A0 (nx2773), .A1 (nx2799)) ;
    mux21 ix2808 (.Y (nx2807), .A0 (nx788), .A1 (nx716), .S0 (nx2849)) ;
    mux21 ix789 (.Y (nx788), .A0 (nx2811), .A1 (nx2813), .S0 (nx726)) ;
    xnor2 ix2812 (.Y (nx2811), .A0 (nx2777), .A1 (nx2793)) ;
    mux21 ix2814 (.Y (nx2813), .A0 (nx780), .A1 (nx732), .S0 (nx2843)) ;
    mux21 ix781 (.Y (nx780), .A0 (nx2817), .A1 (nx2819), .S0 (nx742)) ;
    xnor2 ix2818 (.Y (nx2817), .A0 (nx2781), .A1 (nx2787)) ;
    aoi22 ix2820 (.Y (nx2819), .A0 (nx748), .A1 (T02[2]), .B0 (nx772), .B1 (
          nx750)) ;
    nand02 ix2824 (.Y (nx2823), .A0 (T00[1]), .A1 (T01[0])) ;
    xnor2 ix2826 (.Y (nx2825), .A0 (T00[2]), .A1 (T01[1])) ;
    mux21 ix773 (.Y (nx772), .A0 (nx2829), .A1 (nx2831), .S0 (nx762)) ;
    oai21 ix2830 (.Y (nx2829), .A0 (T01[0]), .A1 (T00[1]), .B0 (nx2823)) ;
    nand02 ix2832 (.Y (nx2831), .A0 (T00[0]), .A1 (T02[0])) ;
    xnor2 ix763 (.Y (nx762), .A0 (T02[1]), .A1 (nx2829)) ;
    xnor2 ix751 (.Y (nx750), .A0 (T02[2]), .A1 (nx2837)) ;
    xnor2 ix2838 (.Y (nx2837), .A0 (nx2823), .A1 (nx2825)) ;
    xnor2 ix743 (.Y (nx742), .A0 (T02[3]), .A1 (nx2817)) ;
    xnor2 ix733 (.Y (nx732), .A0 (nx692), .A1 (nx2789)) ;
    xnor2 ix2844 (.Y (nx2843), .A0 (T02[4]), .A1 (nx732)) ;
    xnor2 ix727 (.Y (nx726), .A0 (T02[5]), .A1 (nx2811)) ;
    xnor2 ix717 (.Y (nx716), .A0 (nx700), .A1 (nx2795)) ;
    xnor2 ix2850 (.Y (nx2849), .A0 (T02[6]), .A1 (nx716)) ;
    xnor2 ix711 (.Y (nx710), .A0 (T02[7]), .A1 (nx2805)) ;
    mux21 ix2856 (.Y (nx2855), .A0 (nx2857), .A1 (nx1156), .S0 (nx1022)) ;
    xnor2 ix2860 (.Y (nx2859), .A0 (T01[7]), .A1 (nx804)) ;
    mux21 ix1157 (.Y (nx1156), .A0 (nx1030), .A1 (nx2865), .S0 (nx1034)) ;
    xnor2 ix1031 (.Y (nx1030), .A0 (nx2807), .A1 (nx710)) ;
    mux21 ix2866 (.Y (nx2865), .A0 (nx2867), .A1 (nx1148), .S0 (nx1046)) ;
    mux21 ix1149 (.Y (nx1148), .A0 (nx1054), .A1 (nx2873), .S0 (nx1058)) ;
    xnor2 ix1055 (.Y (nx1054), .A0 (nx2813), .A1 (nx726)) ;
    mux21 ix2874 (.Y (nx2873), .A0 (nx2875), .A1 (nx1140), .S0 (nx1070)) ;
    mux21 ix1141 (.Y (nx1140), .A0 (nx1078), .A1 (nx2879), .S0 (nx1082)) ;
    xnor2 ix1079 (.Y (nx1078), .A0 (nx2819), .A1 (nx742)) ;
    mux21 ix2880 (.Y (nx2879), .A0 (nx2881), .A1 (nx1132), .S0 (nx1094)) ;
    xnor2 ix2882 (.Y (nx2881), .A0 (nx772), .A1 (nx750)) ;
    mux21 ix1133 (.Y (nx1132), .A0 (nx1102), .A1 (nx2887), .S0 (nx1106)) ;
    xnor2 ix1103 (.Y (nx1102), .A0 (nx2831), .A1 (nx762)) ;
    nor02ii ix2888 (.Y (nx2887), .A0 (nx2889), .A1 (nx2891)) ;
    oai21 ix2890 (.Y (nx2889), .A0 (T02[0]), .A1 (T00[0]), .B0 (nx2831)) ;
    oai21 ix2892 (.Y (nx2891), .A0 (T20[0]), .A1 (T22[0]), .B0 (nx2893)) ;
    nand02 ix2894 (.Y (nx2893), .A0 (T22[0]), .A1 (T20[0])) ;
    xnor2 ix1107 (.Y (nx1106), .A0 (nx1104), .A1 (nx1102)) ;
    xnor2 ix1105 (.Y (nx1104), .A0 (nx2893), .A1 (nx926)) ;
    xnor2 ix927 (.Y (nx926), .A0 (T22[1]), .A1 (nx2901)) ;
    oai21 ix2902 (.Y (nx2901), .A0 (T20[1]), .A1 (T21[0]), .B0 (nx2903)) ;
    nand02 ix2904 (.Y (nx2903), .A0 (T21[0]), .A1 (T20[1])) ;
    xnor2 ix1095 (.Y (nx1094), .A0 (nx2907), .A1 (nx2881)) ;
    xnor2 ix2908 (.Y (nx2907), .A0 (nx936), .A1 (nx914)) ;
    mux21 ix937 (.Y (nx936), .A0 (nx2901), .A1 (nx2893), .S0 (nx926)) ;
    xnor2 ix915 (.Y (nx914), .A0 (T22[2]), .A1 (nx2913)) ;
    xnor2 ix2914 (.Y (nx2913), .A0 (nx2903), .A1 (nx2915)) ;
    xnor2 ix2916 (.Y (nx2915), .A0 (T21[1]), .A1 (T20[2])) ;
    xnor2 ix1083 (.Y (nx1082), .A0 (nx1080), .A1 (nx1078)) ;
    xnor2 ix1081 (.Y (nx1080), .A0 (nx2919), .A1 (nx906)) ;
    aoi22 ix2920 (.Y (nx2919), .A0 (nx912), .A1 (T22[2]), .B0 (nx936), .B1 (
          nx914)) ;
    xnor2 ix907 (.Y (nx906), .A0 (T22[3]), .A1 (nx2925)) ;
    xnor2 ix2926 (.Y (nx2925), .A0 (nx2927), .A1 (nx2933)) ;
    aoi32 ix2928 (.Y (nx2927), .A0 (T21[0]), .A1 (T20[1]), .A2 (nx842), .B0 (
          T20[2]), .B1 (T21[1])) ;
    xnor2 ix2934 (.Y (nx2933), .A0 (T21[2]), .A1 (T20[3])) ;
    xnor2 ix1071 (.Y (nx1070), .A0 (nx1068), .A1 (nx1066)) ;
    xnor2 ix1069 (.Y (nx1068), .A0 (nx944), .A1 (nx2941)) ;
    mux21 ix945 (.Y (nx944), .A0 (nx2925), .A1 (nx2919), .S0 (nx906)) ;
    xnor2 ix2942 (.Y (nx2941), .A0 (T22[4]), .A1 (nx896)) ;
    xnor2 ix897 (.Y (nx896), .A0 (nx856), .A1 (nx2947)) ;
    mux21 ix857 (.Y (nx856), .A0 (nx2927), .A1 (nx2945), .S0 (nx2933)) ;
    inv01 ix2946 (.Y (nx2945), .A (T20[3])) ;
    xnor2 ix2948 (.Y (nx2947), .A0 (T21[3]), .A1 (T20[4])) ;
    xnor2 ix1067 (.Y (nx1066), .A0 (nx780), .A1 (nx2843)) ;
    xnor2 ix1059 (.Y (nx1058), .A0 (nx1056), .A1 (nx1054)) ;
    xnor2 ix1057 (.Y (nx1056), .A0 (nx2955), .A1 (nx890)) ;
    mux21 ix2956 (.Y (nx2955), .A0 (nx944), .A1 (nx896), .S0 (nx2941)) ;
    xnor2 ix891 (.Y (nx890), .A0 (T22[5]), .A1 (nx2959)) ;
    xnor2 ix2960 (.Y (nx2959), .A0 (nx2961), .A1 (nx2963)) ;
    mux21 ix2962 (.Y (nx2961), .A0 (nx856), .A1 (T20[4]), .S0 (nx2947)) ;
    xnor2 ix2964 (.Y (nx2963), .A0 (T21[4]), .A1 (T20[5])) ;
    xnor2 ix1047 (.Y (nx1046), .A0 (nx1044), .A1 (nx1042)) ;
    xnor2 ix1045 (.Y (nx1044), .A0 (nx952), .A1 (nx2971)) ;
    mux21 ix953 (.Y (nx952), .A0 (nx2959), .A1 (nx2955), .S0 (nx890)) ;
    xnor2 ix2972 (.Y (nx2971), .A0 (T22[6]), .A1 (nx880)) ;
    xnor2 ix881 (.Y (nx880), .A0 (nx864), .A1 (nx2979)) ;
    mux21 ix865 (.Y (nx864), .A0 (nx2961), .A1 (nx2977), .S0 (nx2963)) ;
    inv01 ix2978 (.Y (nx2977), .A (T20[5])) ;
    xnor2 ix2980 (.Y (nx2979), .A0 (T21[5]), .A1 (T20[6])) ;
    xnor2 ix1043 (.Y (nx1042), .A0 (nx788), .A1 (nx2849)) ;
    xnor2 ix1035 (.Y (nx1034), .A0 (nx1032), .A1 (nx1030)) ;
    xnor2 ix1033 (.Y (nx1032), .A0 (nx2985), .A1 (nx874)) ;
    mux21 ix2986 (.Y (nx2985), .A0 (nx952), .A1 (nx880), .S0 (nx2971)) ;
    xnor2 ix875 (.Y (nx874), .A0 (T22[7]), .A1 (nx2989)) ;
    xnor2 ix2990 (.Y (nx2989), .A0 (nx2991), .A1 (nx2993)) ;
    mux21 ix2992 (.Y (nx2991), .A0 (nx864), .A1 (T20[6]), .S0 (nx2979)) ;
    xnor2 ix2994 (.Y (nx2993), .A0 (T21[6]), .A1 (T20[7])) ;
    xnor2 ix1023 (.Y (nx1022), .A0 (nx1020), .A1 (nx1014)) ;
    xnor2 ix1021 (.Y (nx1020), .A0 (nx960), .A1 (nx2999)) ;
    mux21 ix961 (.Y (nx960), .A0 (nx2989), .A1 (nx2985), .S0 (nx874)) ;
    xnor2 ix3000 (.Y (nx2999), .A0 (T21[7]), .A1 (nx968)) ;
    mux21 ix969 (.Y (nx968), .A0 (nx2991), .A1 (nx3003), .S0 (nx2993)) ;
    inv01 ix3004 (.Y (nx3003), .A (T20[7])) ;
    xnor2 ix1015 (.Y (nx1014), .A0 (nx796), .A1 (nx2859)) ;
    xnor2 ix1003 (.Y (nx1002), .A0 (nx3009), .A1 (nx3017)) ;
    nor02ii ix3012 (.Y (nx3009), .A0 (nx978), .A1 (nx3015)) ;
    nor02ii ix979 (.Y (nx978), .A0 (nx2999), .A1 (nx960)) ;
    nand02 ix3016 (.Y (nx3015), .A0 (T21[7]), .A1 (nx968)) ;
    nor02ii ix3020 (.Y (nx3017), .A0 (nx814), .A1 (nx2769)) ;
    nor02ii ix815 (.Y (nx814), .A0 (nx2859), .A1 (nx796)) ;
    mux21 ix1263 (.Y (nx1262), .A0 (nx996), .A1 (nx3031), .S0 (nx1002)) ;
    mux21 ix3032 (.Y (nx3031), .A0 (nx3033), .A1 (nx1254), .S0 (nx1022)) ;
    mux21 ix1255 (.Y (nx1254), .A0 (nx1032), .A1 (nx3037), .S0 (nx1034)) ;
    mux21 ix3038 (.Y (nx3037), .A0 (nx3039), .A1 (nx1246), .S0 (nx1046)) ;
    mux21 ix1247 (.Y (nx1246), .A0 (nx1056), .A1 (nx3043), .S0 (nx1058)) ;
    mux21 ix3044 (.Y (nx3043), .A0 (nx3045), .A1 (nx1238), .S0 (nx1070)) ;
    mux21 ix1239 (.Y (nx1238), .A0 (nx1080), .A1 (nx3049), .S0 (nx1082)) ;
    mux21 ix3050 (.Y (nx3049), .A0 (nx2907), .A1 (nx1230), .S0 (nx1094)) ;
    mux21 ix1231 (.Y (nx1230), .A0 (nx1104), .A1 (nx3053), .S0 (nx1106)) ;
    nor02ii ix3054 (.Y (nx3053), .A0 (nx2891), .A1 (nx2889)) ;
    mux21 ix3056 (.Y (nx3055), .A0 (nx3208), .A1 (nx3446), .S0 (nx3295)) ;
    mux21 ix3209 (.Y (nx3208), .A0 (nx3059), .A1 (nx3071), .S0 (nx3715)) ;
    xnor2 ix1285 (.Y (nx1284), .A0 (nx2563), .A1 (nx380)) ;
    xnor2 ix1279 (.Y (nx1278), .A0 (nx2739), .A1 (nx380)) ;
    nand02 ix3068 (.Y (nx3065), .A0 (nx542), .A1 (nx360)) ;
    xnor2 ix1297 (.Y (nx1296), .A0 (nx2855), .A1 (nx1002)) ;
    xnor2 ix1291 (.Y (nx1290), .A0 (nx3031), .A1 (nx1002)) ;
    nand02 ix3078 (.Y (nx3075), .A0 (nx1164), .A1 (nx360)) ;
    mux21 ix3082 (.Y (nx3081), .A0 (nx646), .A1 (nx1598), .S0 (nx3221)) ;
    mux21 ix1599 (.Y (nx1598), .A0 (nx3059), .A1 (nx3085), .S0 (nx3219)) ;
    mux21 ix3086 (.Y (nx3085), .A0 (nx1314), .A1 (nx1582), .S0 (nx3211)) ;
    xnor2 ix3090 (.Y (nx3089), .A0 (nx534), .A1 (nx400)) ;
    xnor2 ix3092 (.Y (nx3091), .A0 (nx632), .A1 (nx400)) ;
    mux21 ix1583 (.Y (nx1582), .A0 (nx3095), .A1 (nx3101), .S0 (nx3203)) ;
    xnor2 ix1337 (.Y (nx1336), .A0 (nx2573), .A1 (nx412)) ;
    xnor2 ix1331 (.Y (nx1330), .A0 (nx2745), .A1 (nx412)) ;
    mux21 ix3102 (.Y (nx3101), .A0 (nx1366), .A1 (nx1566), .S0 (nx3195)) ;
    xnor2 ix3106 (.Y (nx3105), .A0 (nx526), .A1 (nx424)) ;
    xnor2 ix3108 (.Y (nx3107), .A0 (nx624), .A1 (nx424)) ;
    mux21 ix1567 (.Y (nx1566), .A0 (nx3111), .A1 (nx3117), .S0 (nx3187)) ;
    xnor2 ix1389 (.Y (nx1388), .A0 (nx2579), .A1 (nx436)) ;
    xnor2 ix1383 (.Y (nx1382), .A0 (nx2751), .A1 (nx436)) ;
    mux21 ix3118 (.Y (nx3117), .A0 (nx1418), .A1 (nx1550), .S0 (nx3179)) ;
    xnor2 ix3122 (.Y (nx3121), .A0 (nx518), .A1 (nx448)) ;
    xnor2 ix3124 (.Y (nx3123), .A0 (nx616), .A1 (nx448)) ;
    mux21 ix1551 (.Y (nx1550), .A0 (nx3127), .A1 (nx3133), .S0 (nx3171)) ;
    xnor2 ix1441 (.Y (nx1440), .A0 (nx2587), .A1 (nx460)) ;
    xnor2 ix1435 (.Y (nx1434), .A0 (nx2757), .A1 (nx460)) ;
    mux21 ix3134 (.Y (nx3133), .A0 (nx1470), .A1 (nx1534), .S0 (nx3163)) ;
    xnor2 ix3138 (.Y (nx3137), .A0 (nx510), .A1 (nx472)) ;
    xnor2 ix3140 (.Y (nx3139), .A0 (nx608), .A1 (nx472)) ;
    mux21 ix1535 (.Y (nx1534), .A0 (nx3143), .A1 (nx3149), .S0 (nx3155)) ;
    xnor2 ix1493 (.Y (nx1492), .A0 (nx2595), .A1 (nx484)) ;
    xnor2 ix1487 (.Y (nx1486), .A0 (nx2761), .A1 (nx484)) ;
    nand02 ix3150 (.Y (nx3149), .A0 (nx1516), .A1 (nx3153)) ;
    nor02 ix3154 (.Y (nx3153), .A0 (nx3053), .A1 (nx2887)) ;
    xnor2 ix3156 (.Y (nx3155), .A0 (nx3143), .A1 (nx3157)) ;
    xnor2 ix1505 (.Y (nx1504), .A0 (nx2887), .A1 (nx1106)) ;
    xnor2 ix1499 (.Y (nx1498), .A0 (nx3053), .A1 (nx1106)) ;
    xnor2 ix3164 (.Y (nx3163), .A0 (nx1470), .A1 (nx1482)) ;
    xnor2 ix3168 (.Y (nx3167), .A0 (nx1132), .A1 (nx1094)) ;
    xnor2 ix3170 (.Y (nx3169), .A0 (nx1230), .A1 (nx1094)) ;
    xnor2 ix3172 (.Y (nx3171), .A0 (nx3127), .A1 (nx3173)) ;
    xnor2 ix1453 (.Y (nx1452), .A0 (nx2879), .A1 (nx1082)) ;
    xnor2 ix1447 (.Y (nx1446), .A0 (nx3049), .A1 (nx1082)) ;
    xnor2 ix3180 (.Y (nx3179), .A0 (nx1418), .A1 (nx1430)) ;
    xnor2 ix3184 (.Y (nx3183), .A0 (nx1140), .A1 (nx1070)) ;
    xnor2 ix3186 (.Y (nx3185), .A0 (nx1238), .A1 (nx1070)) ;
    xnor2 ix3188 (.Y (nx3187), .A0 (nx3111), .A1 (nx3189)) ;
    xnor2 ix1401 (.Y (nx1400), .A0 (nx2873), .A1 (nx1058)) ;
    xnor2 ix1395 (.Y (nx1394), .A0 (nx3043), .A1 (nx1058)) ;
    xnor2 ix3196 (.Y (nx3195), .A0 (nx1366), .A1 (nx1378)) ;
    xnor2 ix3200 (.Y (nx3199), .A0 (nx1148), .A1 (nx1046)) ;
    xnor2 ix3202 (.Y (nx3201), .A0 (nx1246), .A1 (nx1046)) ;
    xnor2 ix3204 (.Y (nx3203), .A0 (nx3095), .A1 (nx3205)) ;
    xnor2 ix1349 (.Y (nx1348), .A0 (nx2865), .A1 (nx1034)) ;
    xnor2 ix1343 (.Y (nx1342), .A0 (nx3037), .A1 (nx1034)) ;
    xnor2 ix3212 (.Y (nx3211), .A0 (nx1314), .A1 (nx1326)) ;
    xnor2 ix3216 (.Y (nx3215), .A0 (nx1156), .A1 (nx1022)) ;
    xnor2 ix3218 (.Y (nx3217), .A0 (nx1254), .A1 (nx1022)) ;
    xnor2 ix3220 (.Y (nx3219), .A0 (nx3059), .A1 (nx3071)) ;
    xnor2 ix3222 (.Y (nx3221), .A0 (nx646), .A1 (nx1268)) ;
    mux21 ix3447 (.Y (nx3446), .A0 (nx3225), .A1 (nx3227), .S0 (nx3291)) ;
    mux21 ix3226 (.Y (nx3225), .A0 (nx1314), .A1 (nx1326), .S0 (nx3715)) ;
    mux21 ix3228 (.Y (nx3227), .A0 (nx3244), .A1 (nx3430), .S0 (nx3287)) ;
    mux21 ix3245 (.Y (nx3244), .A0 (nx3095), .A1 (nx3205), .S0 (nx3715)) ;
    mux21 ix3431 (.Y (nx3430), .A0 (nx3231), .A1 (nx3233), .S0 (nx3283)) ;
    mux21 ix3232 (.Y (nx3231), .A0 (nx1366), .A1 (nx1378), .S0 (nx3715)) ;
    mux21 ix3234 (.Y (nx3233), .A0 (nx3280), .A1 (nx3414), .S0 (nx3279)) ;
    mux21 ix3281 (.Y (nx3280), .A0 (nx3111), .A1 (nx3189), .S0 (nx3715)) ;
    mux21 ix3415 (.Y (nx3414), .A0 (nx3239), .A1 (nx3241), .S0 (nx3275)) ;
    mux21 ix3240 (.Y (nx3239), .A0 (nx1418), .A1 (nx1430), .S0 (nx3715)) ;
    mux21 ix3242 (.Y (nx3241), .A0 (nx3316), .A1 (nx3398), .S0 (nx3271)) ;
    mux21 ix3317 (.Y (nx3316), .A0 (nx3127), .A1 (nx3173), .S0 (nx3717)) ;
    mux21 ix3399 (.Y (nx3398), .A0 (nx3247), .A1 (nx3249), .S0 (nx3267)) ;
    mux21 ix3248 (.Y (nx3247), .A0 (nx1470), .A1 (nx1482), .S0 (nx3717)) ;
    mux21 ix3250 (.Y (nx3249), .A0 (nx3352), .A1 (nx3382), .S0 (nx3263)) ;
    mux21 ix3353 (.Y (nx3352), .A0 (nx3143), .A1 (nx3157), .S0 (nx3717)) ;
    nor02ii ix3383 (.Y (nx3382), .A0 (nx3378), .A1 (nx3370)) ;
    nor02 ix3258 (.Y (nx3257), .A0 (nx1991), .A1 (nx1813)) ;
    mux21 ix3371 (.Y (nx3370), .A0 (nx3261), .A1 (nx3153), .S0 (nx3717)) ;
    nor02 ix3262 (.Y (nx3261), .A0 (nx2761), .A1 (nx2595)) ;
    xnor2 ix3264 (.Y (nx3263), .A0 (nx3352), .A1 (nx3360)) ;
    xnor2 ix3268 (.Y (nx3267), .A0 (nx3247), .A1 (nx3269)) ;
    xnor2 ix3272 (.Y (nx3271), .A0 (nx3316), .A1 (nx3324)) ;
    xnor2 ix3276 (.Y (nx3275), .A0 (nx3239), .A1 (nx3277)) ;
    xnor2 ix3280 (.Y (nx3279), .A0 (nx3280), .A1 (nx3288)) ;
    xnor2 ix3284 (.Y (nx3283), .A0 (nx3231), .A1 (nx3285)) ;
    xnor2 ix3288 (.Y (nx3287), .A0 (nx3244), .A1 (nx3252)) ;
    xnor2 ix3292 (.Y (nx3291), .A0 (nx3225), .A1 (nx3293)) ;
    xnor2 ix3296 (.Y (nx3295), .A0 (nx3208), .A1 (nx3216)) ;
    xnor2 ix3300 (.Y (nx3299), .A0 (nx2465), .A1 (nx3301)) ;
    nor02 ix3302 (.Y (nx3301), .A0 (nx2852), .A1 (nx2230)) ;
    oai22 ix3893 (.Y (EDGE), .A0 (nx3758), .A1 (nx3547), .B0 (nx3319), .B1 (
          THRESHOLD[10])) ;
    xnor2 ix3759 (.Y (nx3758), .A0 (nx3319), .A1 (THRESHOLD[10])) ;
    xnor2 ix3320 (.Y (nx3319), .A0 (nx3746), .A1 (nx3754)) ;
    nor02 ix3747 (.Y (nx3746), .A0 (nx3323), .A1 (nx3543)) ;
    nand02 ix3324 (.Y (nx3323), .A0 (nx3726), .A1 (nx3734)) ;
    mux21 ix3727 (.Y (nx3726), .A0 (nx3327), .A1 (nx3525), .S0 (nx3537)) ;
    mux21 ix3328 (.Y (nx3327), .A0 (nx3520), .A1 (nx3718), .S0 (nx3530)) ;
    nand02 ix3336 (.Y (nx3335), .A0 (nx3717), .A1 (nx3680)) ;
    mux21 ix3719 (.Y (nx3718), .A0 (nx3357), .A1 (nx3493), .S0 (nx3497)) ;
    mux21 ix3358 (.Y (nx3357), .A0 (nx3576), .A1 (nx3710), .S0 (nx3586)) ;
    mux21 ix3711 (.Y (nx3710), .A0 (nx3381), .A1 (nx3461), .S0 (nx3465)) ;
    mux21 ix3382 (.Y (nx3381), .A0 (nx3632), .A1 (nx3702), .S0 (nx3642)) ;
    mux21 ix3703 (.Y (nx3702), .A0 (nx3405), .A1 (nx3429), .S0 (nx3433)) ;
    aoi221 ix3410 (.Y (nx3409), .A0 (nx3040), .A1 (nx3688), .B0 (nx1444), .B1 (
           nx3686), .C0 (nx3694)) ;
    oai22 ix3695 (.Y (nx3694), .A0 (nx2049), .A1 (nx3719), .B0 (nx3173), .B1 (
          nx3313)) ;
    aoi221 ix3430 (.Y (nx3429), .A0 (nx3014), .A1 (nx3688), .B0 (nx1418), .B1 (
           nx3686), .C0 (nx3658)) ;
    ao22 ix3659 (.Y (nx3658), .A0 (nx3002), .A1 (nx3486), .B0 (nx1430), .B1 (
         nx3478)) ;
    xnor2 ix3434 (.Y (nx3433), .A0 (nx3435), .A1 (nx3429)) ;
    xnor2 ix3643 (.Y (nx3642), .A0 (nx3640), .A1 (nx3441)) ;
    aoi221 ix3442 (.Y (nx3441), .A0 (nx2988), .A1 (nx3688), .B0 (nx1392), .B1 (
           nx3686), .C0 (nx3630)) ;
    oai22 ix3631 (.Y (nx3630), .A0 (nx2033), .A1 (nx3719), .B0 (nx3189), .B1 (
          nx3313)) ;
    aoi221 ix3462 (.Y (nx3461), .A0 (nx2962), .A1 (nx3688), .B0 (nx1366), .B1 (
           nx3686), .C0 (nx3602)) ;
    ao22 ix3603 (.Y (nx3602), .A0 (nx2950), .A1 (nx3486), .B0 (nx1378), .B1 (
         nx3478)) ;
    xnor2 ix3466 (.Y (nx3465), .A0 (nx3467), .A1 (nx3461)) ;
    xnor2 ix3587 (.Y (nx3586), .A0 (nx3584), .A1 (nx3473)) ;
    aoi221 ix3474 (.Y (nx3473), .A0 (nx2936), .A1 (nx3688), .B0 (nx1340), .B1 (
           nx3686), .C0 (nx3574)) ;
    oai22 ix3575 (.Y (nx3574), .A0 (nx2017), .A1 (nx3719), .B0 (nx3205), .B1 (
          nx3313)) ;
    aoi221 ix3494 (.Y (nx3493), .A0 (nx2910), .A1 (nx3472), .B0 (nx1314), .B1 (
           nx3466), .C0 (nx3546)) ;
    ao22 ix3547 (.Y (nx3546), .A0 (nx2898), .A1 (nx3486), .B0 (nx1326), .B1 (
         nx3478)) ;
    xnor2 ix3498 (.Y (nx3497), .A0 (nx3499), .A1 (nx3493)) ;
    xnor2 ix3531 (.Y (nx3530), .A0 (nx3528), .A1 (nx3505)) ;
    aoi221 ix3506 (.Y (nx3505), .A0 (nx2884), .A1 (nx3472), .B0 (nx1288), .B1 (
           nx3466), .C0 (nx3518)) ;
    oai22 ix3519 (.Y (nx3518), .A0 (nx1995), .A1 (nx3719), .B0 (nx3071), .B1 (
          nx3313)) ;
    aoi221 ix3526 (.Y (nx3525), .A0 (nx2230), .A1 (nx3472), .B0 (nx646), .B1 (
           nx3466), .C0 (nx3490)) ;
    xnor2 ix3538 (.Y (nx3537), .A0 (nx3539), .A1 (nx3525)) ;
    nand02 ix3755 (.Y (nx3754), .A0 (nx2465), .A1 (nx3301)) ;
    oai22 ix3877 (.Y (nx3876), .A0 (nx3774), .A1 (nx3555), .B0 (nx3553), .B1 (
          THRESHOLD[8])) ;
    xnor2 ix3775 (.Y (nx3774), .A0 (nx3553), .A1 (THRESHOLD[8])) ;
    xnor2 ix3554 (.Y (nx3553), .A0 (nx3726), .A1 (nx3734)) ;
    oai22 ix3861 (.Y (nx3860), .A0 (nx3782), .A1 (nx3563), .B0 (nx3561), .B1 (
          THRESHOLD[6])) ;
    xnor2 ix3783 (.Y (nx3782), .A0 (nx3561), .A1 (THRESHOLD[6])) ;
    xnor2 ix3562 (.Y (nx3561), .A0 (nx3718), .A1 (nx3530)) ;
    oai22 ix3845 (.Y (nx3844), .A0 (nx3790), .A1 (nx3571), .B0 (nx3569), .B1 (
          THRESHOLD[4])) ;
    xnor2 ix3791 (.Y (nx3790), .A0 (nx3569), .A1 (THRESHOLD[4])) ;
    xnor2 ix3570 (.Y (nx3569), .A0 (nx3710), .A1 (nx3586)) ;
    oai22 ix3829 (.Y (nx3828), .A0 (nx3798), .A1 (nx3579), .B0 (nx3577), .B1 (
          THRESHOLD[2])) ;
    xnor2 ix3799 (.Y (nx3798), .A0 (nx3577), .A1 (THRESHOLD[2])) ;
    xnor2 ix3578 (.Y (nx3577), .A0 (nx3702), .A1 (nx3642)) ;
    xnor2 ix3801 (.Y (nx3800), .A0 (nx3698), .A1 (nx3433)) ;
    nor02 ix3699 (.Y (nx3698), .A0 (nx3407), .A1 (nx3409)) ;
    xnor2 ix3588 (.Y (nx3587), .A0 (nx3407), .A1 (nx3409)) ;
    xnor2 ix3590 (.Y (nx3589), .A0 (nx3800), .A1 (THRESHOLD[1])) ;
    xnor2 ix3795 (.Y (nx3794), .A0 (nx3595), .A1 (THRESHOLD[3])) ;
    xnor2 ix3596 (.Y (nx3595), .A0 (nx3381), .A1 (nx3465)) ;
    xnor2 ix3787 (.Y (nx3786), .A0 (nx3601), .A1 (THRESHOLD[5])) ;
    xnor2 ix3602 (.Y (nx3601), .A0 (nx3357), .A1 (nx3497)) ;
    xnor2 ix3779 (.Y (nx3778), .A0 (nx3607), .A1 (THRESHOLD[7])) ;
    xnor2 ix3608 (.Y (nx3607), .A0 (nx3327), .A1 (nx3537)) ;
    xnor2 ix3767 (.Y (nx3766), .A0 (nx3613), .A1 (THRESHOLD[9])) ;
    xnor2 ix3614 (.Y (nx3613), .A0 (nx3323), .A1 (nx3543)) ;
    aoi21 ix3915 (.Y (DIRECTION[2]), .A0 (nx3313), .A1 (nx3721), .B0 (nx3619)) ;
    oai22 ix3885 (.Y (nx3884), .A0 (nx3766), .A1 (nx3623), .B0 (nx3613), .B1 (
          THRESHOLD[9])) ;
    oai22 ix3869 (.Y (nx3868), .A0 (nx3778), .A1 (nx3627), .B0 (nx3607), .B1 (
          THRESHOLD[7])) ;
    oai22 ix3853 (.Y (nx3852), .A0 (nx3786), .A1 (nx3631), .B0 (nx3601), .B1 (
          THRESHOLD[5])) ;
    oai22 ix3837 (.Y (nx3836), .A0 (nx3794), .A1 (nx3635), .B0 (nx3595), .B1 (
          THRESHOLD[3])) ;
    oai32 ix3821 (.Y (nx3820), .A0 (nx3802), .A1 (nx3587), .A2 (THRESHOLD[0]), .B0 (
          nx3641), .B1 (THRESHOLD[1])) ;
    dffr fsm_inst_reg_state_4 (.Q (O_VALID), .QB (\$dummy [0]), .D (
         fsm_inst_state_3), .CLK (CLOCK), .R (RESET)) ;
    dffr fsm_inst_reg_state_3 (.Q (fsm_inst_state_3), .QB (\$dummy [1]), .D (
         fsm_inst_state_2), .CLK (CLOCK), .R (RESET)) ;
    dffr fsm_inst_reg_state_2 (.Q (fsm_inst_state_2), .QB (\$dummy [2]), .D (
         nx18), .CLK (CLOCK), .R (RESET)) ;
    and02 ix19 (.Y (nx18), .A0 (I_VALID), .A1 (READY)) ;
    dffr fsm_inst_reg_state_1 (.Q (READY), .QB (\$dummy [3]), .D (nx12), .CLK (
         CLOCK), .R (RESET)) ;
    or03 ix13 (.Y (nx12), .A0 (nx8), .A1 (fsm_inst_state_0), .A2 (O_VALID)) ;
    nor02ii ix9 (.Y (nx8), .A0 (I_VALID), .A1 (READY)) ;
    dffs_ni fsm_inst_reg_state_0 (.Q (fsm_inst_state_0), .QB (\$dummy [4]), .D (
            nx1586), .CLK (CLOCK), .S (RESET)) ;
    inv01 ix3548 (.Y (nx3547), .A (nx3884)) ;
    inv01 ix3624 (.Y (nx3623), .A (nx3876)) ;
    inv01 ix3556 (.Y (nx3555), .A (nx3868)) ;
    inv01 ix3628 (.Y (nx3627), .A (nx3860)) ;
    inv01 ix3564 (.Y (nx3563), .A (nx3852)) ;
    inv01 ix3632 (.Y (nx3631), .A (nx3844)) ;
    inv01 ix3572 (.Y (nx3571), .A (nx3836)) ;
    inv01 ix3636 (.Y (nx3635), .A (nx3828)) ;
    inv01 ix3580 (.Y (nx3579), .A (nx3820)) ;
    inv01 ix3803 (.Y (nx3802), .A (nx3589)) ;
    inv01 ix3642 (.Y (nx3641), .A (nx3800)) ;
    inv01 ix3406 (.Y (nx3405), .A (nx3698)) ;
    inv01 ix3633 (.Y (nx3632), .A (nx3441)) ;
    inv01 ix3577 (.Y (nx3576), .A (nx3473)) ;
    inv01 ix3521 (.Y (nx3520), .A (nx3505)) ;
    inv01 ix3314 (.Y (nx3313), .A (nx3478)) ;
    inv01 ix3467 (.Y (nx3466), .A (nx3335)) ;
    inv01 ix3308 (.Y (nx3307), .A (nx3462)) ;
    inv01 ix3101 (.Y (nx3100), .A (nx3257)) ;
    inv01 ix3041 (.Y (nx3040), .A (nx2373)) ;
    inv01 ix2989 (.Y (nx2988), .A (nx2393)) ;
    inv01 ix2937 (.Y (nx2936), .A (nx2415)) ;
    inv01 ix2885 (.Y (nx2884), .A (nx2437)) ;
    inv01 ix2751 (.Y (nx2750), .A (nx2001)) ;
    inv01 ix1984 (.Y (nx1983), .A (nx2652)) ;
    inv01 ix1800 (.Y (nx1799), .A (nx2650)) ;
    inv01 ix1978 (.Y (nx1977), .A (nx2628)) ;
    inv01 ix1792 (.Y (nx1791), .A (nx2626)) ;
    inv01 ix1972 (.Y (nx1971), .A (nx2604)) ;
    inv01 ix1782 (.Y (nx1781), .A (nx2598)) ;
    inv01 ix2581 (.Y (nx2580), .A (nx1943)) ;
    inv01 ix2575 (.Y (nx2574), .A (nx1951)) ;
    inv01 ix2497 (.Y (nx2496), .A (nx1839)) ;
    inv01 ix2427 (.Y (nx2426), .A (nx1841)) ;
    inv01 ix2333 (.Y (nx2332), .A (nx1761)) ;
    inv01 ix2263 (.Y (nx2262), .A (nx1749)) ;
    inv01 ix2129 (.Y (nx2128), .A (nx2115)) ;
    inv01 ix2402 (.Y (nx2401), .A (nx2030)) ;
    inv01 ix2222 (.Y (nx2221), .A (nx2028)) ;
    inv01 ix2424 (.Y (nx2423), .A (nx2006)) ;
    inv01 ix2214 (.Y (nx2213), .A (nx2004)) ;
    inv01 ix2446 (.Y (nx2445), .A (nx1982)) ;
    inv01 ix2204 (.Y (nx2203), .A (nx1976)) ;
    inv01 ix1959 (.Y (nx1958), .A (nx2345)) ;
    inv01 ix1953 (.Y (nx1952), .A (nx2353)) ;
    inv01 ix1875 (.Y (nx1874), .A (nx2241)) ;
    inv01 ix1805 (.Y (nx1804), .A (nx2243)) ;
    inv01 ix1711 (.Y (nx1710), .A (nx2183)) ;
    inv01 ix1641 (.Y (nx1640), .A (nx2177)) ;
    inv01 ix1517 (.Y (nx1516), .A (nx3261)) ;
    inv01 ix1445 (.Y (nx1444), .A (nx3127)) ;
    inv01 ix1393 (.Y (nx1392), .A (nx3111)) ;
    inv01 ix1341 (.Y (nx1340), .A (nx3095)) ;
    inv01 ix1289 (.Y (nx1288), .A (nx3059)) ;
    inv01 ix1167 (.Y (nx1166), .A (nx3075)) ;
    inv01 ix3046 (.Y (nx3045), .A (nx1068)) ;
    inv01 ix2876 (.Y (nx2875), .A (nx1066)) ;
    inv01 ix3040 (.Y (nx3039), .A (nx1044)) ;
    inv01 ix2868 (.Y (nx2867), .A (nx1042)) ;
    inv01 ix3034 (.Y (nx3033), .A (nx1020)) ;
    inv01 ix2858 (.Y (nx2857), .A (nx1014)) ;
    inv01 ix997 (.Y (nx996), .A (nx3009)) ;
    inv01 ix991 (.Y (nx990), .A (nx3017)) ;
    inv01 ix913 (.Y (nx912), .A (nx2913)) ;
    inv01 ix843 (.Y (nx842), .A (nx2915)) ;
    inv01 ix749 (.Y (nx748), .A (nx2837)) ;
    inv01 ix679 (.Y (nx678), .A (nx2825)) ;
    inv01 ix545 (.Y (nx544), .A (nx3065)) ;
    inv01 ix2754 (.Y (nx2753), .A (nx446)) ;
    inv01 ix2582 (.Y (nx2581), .A (nx444)) ;
    inv01 ix2748 (.Y (nx2747), .A (nx422)) ;
    inv01 ix2576 (.Y (nx2575), .A (nx420)) ;
    inv01 ix2742 (.Y (nx2741), .A (nx398)) ;
    inv01 ix2566 (.Y (nx2565), .A (nx392)) ;
    inv01 ix375 (.Y (nx374), .A (nx2717)) ;
    inv01 ix369 (.Y (nx368), .A (nx2725)) ;
    inv01 ix291 (.Y (nx290), .A (nx2621)) ;
    inv01 ix221 (.Y (nx220), .A (nx2623)) ;
    inv01 ix127 (.Y (nx126), .A (nx2545)) ;
    inv01 ix57 (.Y (nx56), .A (nx2533)) ;
    inv01 ix3620 (.Y (nx3619), .A (EDGE)) ;
    inv01 ix3679 (.Y (nx3680), .A (nx3735)) ;
    inv01 ix3685 (.Y (nx3686), .A (nx3335)) ;
    inv01 ix3689 (.Y (nx3690), .A (nx1957)) ;
    buf02 ix3714 (.Y (nx3715), .A (nx3081)) ;
    buf02 ix3716 (.Y (nx3717), .A (nx3081)) ;
    inv01 ix3718 (.Y (nx3719), .A (nx3486)) ;
    inv01 ix3720 (.Y (nx3721), .A (nx3486)) ;
    and02 ix3473 (.Y (nx3472), .A0 (nx3739), .A1 (nx3735)) ;
    nor02ii ix2853 (.Y (nx2852), .A0 (nx2846), .A1 (nx2001)) ;
    mux21 ix1996 (.Y (nx1995), .A0 (nx2862), .A1 (nx2868), .S0 (nx3733)) ;
    mux21 ix2899 (.Y (nx2898), .A0 (nx2013), .A1 (nx2011), .S0 (nx3733)) ;
    mux21 ix2018 (.Y (nx2017), .A0 (nx2914), .A1 (nx2920), .S0 (nx3733)) ;
    mux21 ix2951 (.Y (nx2950), .A0 (nx2029), .A1 (nx2027), .S0 (nx3733)) ;
    mux21 ix2034 (.Y (nx2033), .A0 (nx2966), .A1 (nx2972), .S0 (nx3733)) ;
    mux21 ix3003 (.Y (nx3002), .A0 (nx2045), .A1 (nx2043), .S0 (nx2750)) ;
    mux21 ix2050 (.Y (nx2049), .A0 (nx3018), .A1 (nx3024), .S0 (nx2750)) ;
    mux21 ix3055 (.Y (nx3054), .A0 (nx2061), .A1 (nx2059), .S0 (nx2750)) ;
    mux21 ix2066 (.Y (nx2065), .A0 (nx3070), .A1 (nx3076), .S0 (nx2750)) ;
    mux21 ix2092 (.Y (nx2091), .A0 (nx3082), .A1 (nx3088), .S0 (nx3731)) ;
    mux21 ix3067 (.Y (nx3066), .A0 (nx2367), .A1 (nx2365), .S0 (nx3731)) ;
    mux21 ix2374 (.Y (nx2373), .A0 (nx3030), .A1 (nx3036), .S0 (nx3731)) ;
    mux21 ix3015 (.Y (nx3014), .A0 (nx2387), .A1 (nx2385), .S0 (nx3731)) ;
    mux21 ix2394 (.Y (nx2393), .A0 (nx2978), .A1 (nx2984), .S0 (nx3731)) ;
    mux21 ix2963 (.Y (nx2962), .A0 (nx2409), .A1 (nx2407), .S0 (nx3731)) ;
    mux21 ix2416 (.Y (nx2415), .A0 (nx2926), .A1 (nx2932), .S0 (nx2128)) ;
    mux21 ix2911 (.Y (nx2910), .A0 (nx2431), .A1 (nx2429), .S0 (nx2128)) ;
    mux21 ix2438 (.Y (nx2437), .A0 (nx2874), .A1 (nx2880), .S0 (nx2128)) ;
    nor02ii ix2231 (.Y (nx2230), .A0 (nx2224), .A1 (nx2115)) ;
    nor02ii ix647 (.Y (nx646), .A0 (nx640), .A1 (nx3065)) ;
    nor02ii ix1269 (.Y (nx1268), .A0 (nx1262), .A1 (nx3075)) ;
    mux21 ix3060 (.Y (nx3059), .A0 (nx1278), .A1 (nx1284), .S0 (nx3727)) ;
    mux21 ix3072 (.Y (nx3071), .A0 (nx1290), .A1 (nx1296), .S0 (nx3729)) ;
    mux21 ix1315 (.Y (nx1314), .A0 (nx3091), .A1 (nx3089), .S0 (nx3727)) ;
    mux21 ix3096 (.Y (nx3095), .A0 (nx1330), .A1 (nx1336), .S0 (nx3727)) ;
    mux21 ix1367 (.Y (nx1366), .A0 (nx3107), .A1 (nx3105), .S0 (nx3727)) ;
    mux21 ix3112 (.Y (nx3111), .A0 (nx1382), .A1 (nx1388), .S0 (nx3727)) ;
    mux21 ix1419 (.Y (nx1418), .A0 (nx3123), .A1 (nx3121), .S0 (nx3727)) ;
    mux21 ix3128 (.Y (nx3127), .A0 (nx1434), .A1 (nx1440), .S0 (nx544)) ;
    mux21 ix1471 (.Y (nx1470), .A0 (nx3139), .A1 (nx3137), .S0 (nx544)) ;
    mux21 ix3144 (.Y (nx3143), .A0 (nx1486), .A1 (nx1492), .S0 (nx544)) ;
    mux21 ix3158 (.Y (nx3157), .A0 (nx1498), .A1 (nx1504), .S0 (nx3729)) ;
    mux21 ix1483 (.Y (nx1482), .A0 (nx3169), .A1 (nx3167), .S0 (nx3729)) ;
    mux21 ix3174 (.Y (nx3173), .A0 (nx1446), .A1 (nx1452), .S0 (nx3729)) ;
    mux21 ix1431 (.Y (nx1430), .A0 (nx3185), .A1 (nx3183), .S0 (nx3729)) ;
    mux21 ix3190 (.Y (nx3189), .A0 (nx1394), .A1 (nx1400), .S0 (nx1166)) ;
    mux21 ix1379 (.Y (nx1378), .A0 (nx3201), .A1 (nx3199), .S0 (nx1166)) ;
    mux21 ix3206 (.Y (nx3205), .A0 (nx1342), .A1 (nx1348), .S0 (nx1166)) ;
    mux21 ix1327 (.Y (nx1326), .A0 (nx3217), .A1 (nx3215), .S0 (nx1166)) ;
    mux21 ix3379 (.Y (nx3378), .A0 (nx2075), .A1 (nx3257), .S0 (nx3739)) ;
    mux21 ix3361 (.Y (nx3360), .A0 (nx2091), .A1 (nx2065), .S0 (nx3739)) ;
    mux21 ix3270 (.Y (nx3269), .A0 (nx3066), .A1 (nx3054), .S0 (nx3739)) ;
    mux21 ix3325 (.Y (nx3324), .A0 (nx2373), .A1 (nx2049), .S0 (nx3739)) ;
    mux21 ix3278 (.Y (nx3277), .A0 (nx3014), .A1 (nx3002), .S0 (nx3739)) ;
    mux21 ix3289 (.Y (nx3288), .A0 (nx2393), .A1 (nx2033), .S0 (nx3741)) ;
    mux21 ix3286 (.Y (nx3285), .A0 (nx2962), .A1 (nx2950), .S0 (nx3741)) ;
    mux21 ix3253 (.Y (nx3252), .A0 (nx2415), .A1 (nx2017), .S0 (nx3741)) ;
    mux21 ix3294 (.Y (nx3293), .A0 (nx2910), .A1 (nx2898), .S0 (nx3741)) ;
    mux21 ix3217 (.Y (nx3216), .A0 (nx2437), .A1 (nx1995), .S0 (nx3741)) ;
    ao22 ix3905 (.Y (nx3904), .A0 (nx2128), .A1 (nx3486), .B0 (nx544), .B1 (
         nx3478)) ;
    nor02 ix3312 (.Y (nx3486), .A0 (nx3741), .A1 (nx3462)) ;
    nor02ii ix3479 (.Y (nx3478), .A0 (nx3717), .A1 (nx3462)) ;
    mux21 ix3408 (.Y (nx3407), .A0 (nx3370), .A1 (nx3378), .S0 (nx3735)) ;
    mux21 ix3436 (.Y (nx3435), .A0 (nx3352), .A1 (nx3360), .S0 (nx3735)) ;
    mux21 ix3641 (.Y (nx3640), .A0 (nx3247), .A1 (nx3269), .S0 (nx3735)) ;
    mux21 ix3468 (.Y (nx3467), .A0 (nx3316), .A1 (nx3324), .S0 (nx3735)) ;
    mux21 ix3585 (.Y (nx3584), .A0 (nx3239), .A1 (nx3277), .S0 (nx3737)) ;
    mux21 ix3500 (.Y (nx3499), .A0 (nx3280), .A1 (nx3288), .S0 (nx3737)) ;
    mux21 ix3529 (.Y (nx3528), .A0 (nx3231), .A1 (nx3285), .S0 (nx3737)) ;
    ao22 ix3491 (.Y (nx3490), .A0 (nx2852), .A1 (nx3486), .B0 (nx1268), .B1 (
         nx3478)) ;
    mux21 ix3540 (.Y (nx3539), .A0 (nx3244), .A1 (nx3252), .S0 (nx3737)) ;
    mux21 ix3735 (.Y (nx3734), .A0 (nx3225), .A1 (nx3293), .S0 (nx3737)) ;
    mux21 ix3544 (.Y (nx3543), .A0 (nx3208), .A1 (nx3216), .S0 (nx3737)) ;
    nor02ii ix3911 (.Y (DIRECTION[1]), .A0 (nx3307), .A1 (EDGE)) ;
    and02 ix3687 (.Y (nx3688), .A0 (nx3690), .A1 (nx3307)) ;
    inv01 ix3726 (.Y (nx3727), .A (nx3065)) ;
    inv01 ix3728 (.Y (nx3729), .A (nx3075)) ;
    inv01 ix3730 (.Y (nx3731), .A (nx2115)) ;
    inv01 ix3732 (.Y (nx3733), .A (nx2001)) ;
    inv01 ix3734 (.Y (nx3735), .A (nx3462)) ;
    inv01 ix3736 (.Y (nx3737), .A (nx3462)) ;
    inv01 ix3738 (.Y (nx3739), .A (nx1957)) ;
    inv01 ix3740 (.Y (nx3741), .A (nx1957)) ;
endmodule

