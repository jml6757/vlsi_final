  X �     �      mentor.db  >A�7KƧ�9D�/��ZP �     �      via4        ,���<���<  	����<  	�  	����<  	����<���<      !    ,���<���<  	����<  	�  	����<  	����<���<           ,���$���$  ����$  �  ����$  ����$���$     �     �      via3    >    ,���<���<  	����<  	�  	����<  	����<���<          ,���<���<  	����<  	�  	����<  	����<���<          ,���$���$  ����$  �  ����$  ����$���$     �     �      via2    3    ,���<���<  	����<  	�  	����<  	����<���<      >    ,���<���<  	����<  	�  	����<  	����<���<      =    ,���$���$  ����$  �  ����$  ����$���$     �    	 %�    	 & via     1    ,���<���<  	����<  	�  	����<  	����<���<      3    ,���<���<  	����<  	�  	����<  	����<���<      2    ,���$���$  ����$  �  ����$  ����$���$     �   
   '� 	   1  
oai32     0    ,  �\  [�  ��  [�  ��  c�  �\  c�  �\  [�      0    ,  �\  s<  ��  s<  ��  {  �\  {  �\  s<      1    ,  �D  W�  ��  W�  ��  ~�  �D  ~�  �D  W� +  ,1       .    ,  ��  L,  ��  L,  ��  U�  ��  U�  ��  L, +  ,3       .    ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� +  ,4       .    ,  ��  U�  ��  U�  ��  ��  ��  ��  ��  U�      0    ,  �  [�  �L  [�  �L  c�  �  c�  �  [�      0    ,  �  s<  �L  s<  �L  {  �  {  �  s<      1    ,  �  W�  �d  W�  �d  ~�  �  ~�  �  W� +  ,5       .    ,  �|  L,  ��  L,  ��  U�  �|  U�  �|  L, +  ,6       .    ,  �|  ��  ��  ��  ��  ��  �|  ��  �|  �� +  ,7       .    ,  �|  U�  ��  U�  ��  ��  �|  ��  �|  U�      0    ,  ��  [�  {  [�  {  c�  ��  c�  ��  [�      0    ,  ��  s<  {  s<  {  {  ��  {  ��  s<      1    ,  ��  W�  w$  W�  w$  ~�  ��  ~�  ��  W� +  ,8       .    ,  s<  L,  kl  L,  kl  U�  s<  U�  s<  L, +  ,9       .    ,  s<  ��  kl  ��  kl  ��  s<  ��  s<  �� +  ,10      .    ,  s<  U�  kl  U�  kl  ��  s<  ��  s<  U�      0    ,  c�  [�  [�  [�  [�  c�  c�  c�  c�  [�      0    ,  c�  s<  [�  s<  [�  {  c�  {  c�  s<      1    ,  g�  W�  W�  W�  W�  ~�  g�  ~�  g�  W� +  ,11      .    ,  S�  L,  L,  L,  L,  U�  S�  U�  S�  L, +  ,12      .    ,  S�  ��  L,  ��  L,  ��  S�  ��  S�  �� +  ,13      .    ,  S�  U�  L,  U�  L,  ��  S�  ��  S�  U�      0    ,  D\  [�  <�  [�  <�  c�  D\  c�  D\  [�      0    ,  D\  s<  <�  s<  <�  {  D\  {  D\  s<      1    ,  HD  W�  8�  W�  8�  ~�  HD  ~�  HD  W� +  ,14      .    ,  4�  L,  ,�  L,  ,�  U�  4�  U�  4�  L, +  ,15      .    ,  4�  ��  ,�  ��  ,�  ��  4�  ��  4�  �� +  ,16      .    ,  4�  U�  ,�  U�  ,�  ��  4�  ��  4�  U�      0    ,  %  [�  L  [�  L  c�  %  c�  %  [�      0    ,  %  s<  L  s<  L  {  %  {  %  s<      +    ,  �8  U�  ��  U�  ��  ��  �8  ��  �8  U� +  ,2       1    ,  )  W�  d  W�  d  ~�  )  ~�  )  W� +  ,17      +    ,  �8  U�  p  U�  p  ��  �8  ��  �8  U�      )    ,  ި  >�      >�      �X  ި  �X  ި  >� +  ,19      -    ,  �  N   �  N   �  ��  �  ��  �  N       +    ,  ,�  U�  p  U�  p  ��  ,�  ��  ,�  U� +  ,18      0    ,  ��  ��  ��  ��  �� �  �� �  ��  ��      0    ,  �� L  �� L  ��   ��   �� L      0    ,  �� .�  �� .�  �� 6�  �� 6�  �� .�      0    ,  �� F,  �� F,  �� M�  �� M�  �� F,      0    ,  �� ]�  �� ]�  �� el  �� el  �� ]�      1    ,  �h  ��  ��  ��  �� iT  �h iT  �h  �� +  ,1       .    ,  ��  �<  �  �<  �  �   ��  �   ��  �< +  ,3       .    ,  �� kH  � kH  � u  �� u  �� kH +  ,4       .    ,  ��  �   �  �   � kH  �� kH  ��  �       .    ,  �p  �<  ��  �<  ��  �   �p  �   �p  �< +  ,5       .    ,  �p kH  �� kH  �� u  �p u  �p kH +  ,6       .    ,  �p  �   ��  �   �� kH  �p kH  �p  �       0    ,  ��  ��  {  ��  { �  �� �  ��  ��      0    ,  �� L  { L  {   ��   �� L      0    ,  �� .�  { .�  { 6�  �� 6�  �� .�      0    ,  �� F,  { F,  { M�  �� M�  �� F,      0    ,  �� ]�  { ]�  { el  �� el  �� ]�      0    ,  �� u  { u  { |�  �� |�  �� u      0    ,  �� �|  { �|  { �L  �� �L  �� �|      1    ,  ��  ��  w$  ��  w$ �4  �� �4  ��  �� +  ,7       .    ,  s<  �<  kl  �<  kl  �   s<  �   s<  �< +  ,8       .    ,  s< ��  kl ��  kl ��  s< ��  s< �� +  ,9       .    ,  s<  �   kl  �   kl ��  s< ��  s<  �       .    ,  [�  �<  S�  �<  S�  �   [�  �   [�  �< +  ,10      .    ,  [� ��  S� ��  S� ��  [� ��  [� �� +  ,11      .    ,  [�  �   S�  �   S� ��  [� ��  [�  �       .    ,  D\  �<  <�  �<  <�  �   D\  �   D\  �< +  ,12      .    ,  D\ ��  <� ��  <� ��  D\ ��  D\ �� +  ,13      .    ,  D\  �   <�  �   <� ��  D\ ��  D\  �       0    ,  4� �  ,� �  ,� |  4� |  4� �      0    ,  4�   ,�   ,� &�  4� &�  4�       0    ,  4� 6�  ,� 6�  ,� >\  4� >\  4� 6�      0    ,  4� M�  ,� M�  ,� U�  4� U�  4� M�      0    ,  4� el  ,� el  ,� m<  4� m<  4� el      0    ,  4� |�  ,� |�  ,� ��  4� ��  4� |�      0    ,  4� �L  ,� �L  ,� �  4� �  4� �L      +    ,  �\  �   ��  �   �� kH  �\ kH  �\  �  +  ,2       1    ,  8� �  ) �  ) �  8� �  8� � +  ,14      +    \  ,�  �   ,� �  ' �  ' ��  �� ��  �� �(  �� �(  �� kH  �\ kH  �\  �   ,�  �       *    \  |  �  |  �`  �  �`  � �h  �L �h  �L ��  �( ��  �( ��  �� ��  ��  �  |  � +  ,16      ,    \  %  �0  %  �   @  �   @ ��  �� ��  �� ��  �� ��  �� s  �, s  �,  �0  %  �0      +    <  ,�  �   ,� �  ' �  ' ��  <� ��  <�  �   ,�  �  +  ,15   
  via    ��  �P   
  via    <�  �P   
  via    �  �P   
  via    _�  �P   
  via    �,  �P   
  via    d  �P      3    ,  2�  ��  FP  ��  FP  �  2�  �  2�  ��      3    ,  �h  ��  ��  ��  ��  �  �h  �  �h  ��      3    ,  y  ��  ��  ��  ��  �  y  �  y  ��      3    ,  �@  ��  ��  ��  ��  �  �@  �  �@  ��      3    ,  U�  ��  ix  ��  ix  �  U�  �  U�  ��      3    ,  �  ��  #(  ��  #(  �  �  �  �  ��      1    ,          ި      ި  '      '              1    ,     ��  ި ��  ި ��     ��     ��      �    ,          ި      ި ��     ��           	   .      � $  ��  �<  ��  ��  �(  ��  �(  �      .    ,  ix  ��  kl  ��  kl  �  ix  �  ix  ��   	   .      �   ��  ��  �P  ��  �P  ��      .    ,  U�  ��  ix  ��  ix  �  U�  �  U�  ��      .    ,  2�  ��  FP  ��  FP  �  2�  �  2�  ��   	   .      �   �  �T  �P  �T  �P  �      .    ,  �@  ��  ��  ��  ��  �  �@  �  �@  ��   	   .      �   4�  ��  @  ��  @  ��      .    ,  �h  ��  ��  ��  ��  �  �h  �  �h  ��      .    ,  �  ��  #(  ��  #(  �  �  �  �  ��   	   .      �   D\  �0  @  �0  @  �   	   .      �   oT  �<  oT  ��   	   .      � $  Bh  ��  Bh  �  P  �  P  ��   	   .      � $  �(  ��  �(  ��  ��  ��  ��  ��   	   .      � $  W�  �<  W�  ި  Bh  ި  Bh  �      /    ,  8�  �h  @t  �h  @t  �8  8�  �8  8�  �h      /    ,  �  �h  ��  �h  ��  �8  �  �8  �  �h      /    ,  �D  �h  �  �h  �  �8  �D  �8  �D  �h      /    ,  [�  �h  c�  �h  c�  �8  [�  �8  [�  �h      /    ,  |  �h  L  �h  L  �8  |  �8  |  �h      -    ,  � ��  �� ��  �� ��  � ��  � ��      -    ,  � s  �, s  �, ��  � ��  � s      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      ,    ,  ��  *�  ��  *�  ��  N   ��  N   ��  *�      0    ,  0�  |  8�  |  8�  L  0�  L  0�  |      0    ,  HD  |  P  |  P  L  HD  L  HD  |      0    ,  w$  |  ~�  |  ~�  L  w$  L  w$  |      0    ,  _�  |  g�  |  g�  L  _�  L  _�  |      0    ,  �  |  ��  |  ��  L  �  L  �  |      0    ,  ��  |  �d  |  �d  L  ��  L  ��  |      0    ,  �t  |  �D  |  �D  L  �t  L  �t  |      0    ,  d  |  !4  |  !4  L  d  L  d  |      0    ,  �� �t  �d �t  �d �D  �� �D  �� �t      0    ,  w$ �t  ~� �t  ~� �D  w$ �D  w$ �t      0    ,  _� �t  g� �t  g� �D  _� �D  _� �t      0    ,  HD �t  P �t  P �D  HD �D  HD �t      0    ,  0� �t  8� �t  8� �D  0� �D  0� �t      0    ,  d �t  !4 �t  !4 �D  d �D  d �t      0    ,  � �t  �� �t  �� �D  � �D  � �t      0    ,  �t �t  �D �t  �D �D  �t �D  �t �t      0    ,  �� ��  �� ��  �� ��  �� ��  �� ��      0    ,  �� �  �� �  �� ��  �� ��  �� �      0    ,  �L  8�  �  8�  �  @t  �L  @t  �L  8�      1    ,  �\  ��  ��  ��  ��  �   �\  �   �\  ��      1    ,  �4  ��  ��  ��  ��  �   �4  �   �4  ��   	   1      �   ~�  �  ~�  ��      1    ,  �� iT  �h iT  �h z�  �� z�  �� iT   	   1      � $  �t  ~�  �t  ��  ~�  ��  ~�  ~�      1    ,  W�  ��  g�  ��  g�  �   W�  �   W�  ��      1    ,  �  ��  !4  ��  !4  �   �  �   �  ��      1    ,  ) �  6� �  6� ��  ) ��  ) �   	   1      � $  _�  ~�  _�  ��  !4  ��  !4  ~�   	   1      � $  ~�  W�  ~�  >�  @t  >�  @t  W�      1    ,  4�  ��  D\  ��  D\  �   4�  �   4�  ��   	   1      � $  ~�  ��  ~�  ��  _�  ��  _�  �d      1    ,  �� z�  �h z�  �h ��  �� ��  �� z�      1    ,  �X  D\  �  D\  �  W�  �X  W�  �X  D\      1    ,  �d  '  �  '  �  D\  �d  D\  �d  '      +    ,  �  �  �   �  �   #(  �  #(  �  �      +    ,  � ��  �  ��  �  �   � �   � ��      +    ,  ' ��  8� ��  8� ��  ' ��  ' ��      +    ,  �� x�  �\ x�  �\ ��  �� ��  �� x�      +    ,  �� kH  �\ kH  �\ x�  �� x�  �� kH      +    ,  �d  FP  �  FP  �  U�  �d  U�  �d  FP      +    ,  �p  #(  ��  #(  ��  FP  �p  FP  �p  #(      *    ,      �  ި  �  ި ��     ��      �      )    ,          ި      ި  �X      �X                      oT  � GND  +  ,1               oT �8 VDD  +  ,1               ��  �P Y  +  ,1               _�  �P A2 +  ,1               �  �P B1 +  ,1               <�  �P A1 +  ,1               d  �P A0 +  ,1               �,  �P B0 +  ,1               oT  � GND               oT �8 VDD               ��  �P Y               _�  �P A2              �  �P B1              <�  �P A1              d  �P A0              �,  �P B0     �     � 	   / - 
buf02     +    ,  kl X  U� X  U� @P  kl @P  kl X +  ,2       0    ,  e� 4  ]� 4  ]� #  e� #  e� 4      0    ,  e� 2�  ]� 2�  ]� :t  e� :t  e� 2�      1    ,  ix L  Y� L  Y� >\  ix >\  ix L +  ,1       .    ,  U� �  N  �  N  X  U� X  U� � +  ,3       .    ,  U� @P  N  @P  N  J  U� J  U� @P +  ,4       .    ,  U� X  N  X  N  @P  U� @P  U� X      0    ,  D\ .�  <� .�  <� 6�  D\ 6�  D\ .�      0    ,  D\ F,  <� F,  <� M�  D\ M�  D\ F,      0    ,  D\ ]�  <� ]�  <� el  D\ el  D\ ]�      1    ,  HD *�  8� *�  8� iT  HD iT  HD *� +  ,5       .    ,  4� �  ,� �  ,� X  4� X  4� � +  ,6       .    ,  4� kH  ,� kH  ,� u  4� u  4� kH +  ,7       .    ,  4� X  ,� X  ,� kH  4� kH  4� X      0    ,  % 4  L 4  L #  % #  % 4      0    ,  % 2�  L 2�  L :t  % :t  % 2�      0    ,  % J  L J  L Q�  % Q�  % J      1    ,  ) L  d L  d U�  ) U�  ) L +  ,8       +    L  p X  p W�  L W�  L kH  J8 kH  J8 @P  kl @P  kl X  p X      *    L      ��     o0  � o0  � ��  a� ��  a� W�  �� W�  ��  ��      �� +  ,10      ,    L  � �  � _�  | _�  | s  R s  R H   s< H   s< �  � �      +    <  p X  p W�  L W�  L kH  ,� kH  ,� X  p X +  ,9       +    ,  p  a�  ,�  a�  ,�  ��  p  ��  p  a� +  ,2       0    ,  L  g�  %  g�  %  oT  L  oT  L  g�      0    ,  L  ~�  %  ~�  %  ��  L  ��  L  ~�      1    ,  d  c�  )  c�  )  ��  d  ��  d  c� +  ,1       .    ,  ,�  W�  4�  W�  4�  a�  ,�  a�  ,�  W� +  ,3       .    ,  ,�  ��  4�  ��  4�  �d  ,�  �d  ,�  �� +  ,4       .    ,  ,�  a�  4�  a�  4�  ��  ,�  ��  ,�  a�      0    ,  <�  g�  D\  g�  D\  oT  <�  oT  <�  g�      0    ,  <�  ~�  D\  ~�  D\  ��  <�  ��  <�  ~�      1    ,  8�  c�  HD  c�  HD  ��  8�  ��  8�  c� +  ,5       .    ,  N   oT  U�  oT  U�  y  N   y  N   oT +  ,6       .    ,  N   ��  U�  ��  U�  �d  N   �d  N   �� +  ,7       .    ,  N   y  U�  y  U�  ��  N   ��  N   y      0    ,  ]�  ~�  e�  ~�  e�  ��  ]�  ��  ]�  ~�      1    ,  Y�  {  ix  {  ix  ��  Y�  ��  Y�  { +  ,8       +    <  J8  a�  J8  y  kl  y  kl  ��  p  ��  p  a�  J8  a�      )    <  a�  J8  a�  a�  ��  a�  ��  �      �      J8  a�  J8 +  ,10      -    <  R  Y�  R  qH  s<  qH  s<  �p  �  �p  �  Y�  R  Y�      +    ,  U�  y  kl  y  kl  ��  U�  ��  U�  y +  ,9    
  via     BZ         L,  �   
  via    L  �      3    ,  Bh  �P  U�  �P  U�  ��  Bh  ��  Bh  �P      3    ,  �  �P  '  �P  '  ��  �  ��  �  �P      1    ,     ��  �� ��  �� ��     ��     ��      1    ,          ��      ��  '      '              0    ,  0�  |  8�  |  8�  L  0�  L  0�  |      0    ,  HD  |  P  |  P  L  HD  L  HD  |      0    ,  _�  |  g�  |  g�  L  _�  L  _�  |      0    ,  d  |  !4  |  !4  L  d  L  d  |      0    ,  d �t  !4 �t  !4 �D  d �D  d �t      0    ,  0� �t  8� �t  8� �D  0� �D  0� �t      0    ,  HD �t  P �t  P �D  HD �D  HD �t      0    ,  _� �t  g� �t  g� �D  _� �D  _� �t      0    ,  <�  D\  D\  D\  D\  L,  <�  L,  <�  D\      0    ,  <�  ,�  D\  ,�  D\  4�  <�  4�  <�  ,�      0    ,  <� ��  D\ ��  D\ ��  <� ��  <� ��      0    ,  <� �4  D\ �4  D\ �  <� �  <� �4      1    ,  D\  �D  S�  �D  S�  ��  D\  ��  D\  �D   	   1      �   g�  ~�  g� #   	   1      �   @ L  @  ��   	   1      �   @  �P  @  ��      1    ,  :� iT  HD iT  HD |�  :� |�  :� iT      1    ,  8� |�  HD |�  HD ��  8� ��  8� |�      1    ,  0�  �   @t  �   @t 	�  0� 	�  0�  �    	   1      �   @t �  a� �      1    ,  8�  '  HD  '  HD  P  8�  P  8�  '      1    ,  :�  P  HD  P  HD  c�  :�  c�  :�  P      +    ,  �  �  m`  �  m`  #(  �  #(  �  �      +    ,  � ��  m` ��  m` �   � �   � ��      +    ,  6�  #(  J8  #(  J8  R  6�  R  6�  #(      +    ,  8�  R  J8  R  J8  a�  8�  a�  8�  R      +    ,  6� z�  J8 z�  J8 ��  6� ��  6� z�      +    ,  8� kH  J8 kH  J8 z�  8� z�  8� kH      -    ,  � ��  u0 ��  u0 ��  � ��  � ��      -    ,  .� s  R s  R ��  .� ��  .� s      ,    ,  �  �  u0  �  u0  *�  �  *�  �  �      ,    ,  .�  *�  R  *�  R  Y�  .�  Y�  .�  *�      )    ,          ��      ��  �      �              *    ,      ��  ��  ��  �� ��     ��      ��      /    ,  HD  �,  P  �,  P  ��  HD  ��  HD  �,      /    ,  4�  ��  <�  ��  <� �  4� �  4�  ��      .    ,  Bh  �P  U�  �P  U�  ��  Bh  ��  Bh  �P      .    ,  .�  �  Bh  �  Bh �  .� �  .�  �   	   .      �   R �  R  ��   	   .      �   0� �  0�  �d   	   .      �   R  �d  R  �P              An  � GND  +  ,1               An �8 VDD  +  ,1               L  � Y  +  ,1               L,  � A  +  ,1       �    ,          ��      �� ��     ��                      An  � GND               An �8 VDD               L  � Y               L,  � A      �   	 1 (� 	   /  
aoi21     +    ,  �� (�  s< (�  s< kH  �� kH  �� (� +  ,2       0    ,  �� .�  { .�  { 6�  �� 6�  �� .�      0    ,  �� F,  { F,  { M�  �� M�  �� F,      0    ,  �� ]�  { ]�  { el  �� el  �� ]�      1    ,  �� *�  w$ *�  w$ iT  �� iT  �� *� +  ,1       .    ,  s<   kl   kl (�  s< (�  s<  +  ,3       .    ,  s< kH  kl kH  kl u  s< u  s< kH +  ,4       .    ,  s< (�  kl (�  kl kH  s< kH  s< (�      0    ,  c� .�  [� .�  [� 6�  c� 6�  c� .�      0    ,  c� F,  [� F,  [� M�  c� M�  c� F,      0    ,  c� ]�  [� ]�  [� el  c� el  c� ]�      1    ,  g� *�  W� *�  W� iT  g� iT  g� *� +  ,5       .    ,  S�   L,   L, (�  S� (�  S�  +  ,6       .    ,  S� kH  L, kH  L, u  S� u  S� kH +  ,7       .    ,  S� (�  L, (�  L, kH  S� kH  S� (�      0    ,  D\ .�  <� .�  <� 6�  D\ 6�  D\ .�      0    ,  D\ F,  <� F,  <� M�  D\ M�  D\ F,      0    ,  D\ ]�  <� ]�  <� el  D\ el  D\ ]�      1    ,  HD *�  8� *�  8� iT  HD iT  HD *� +  ,8       .    ,  4�   ,�   ,� (�  4� (�  4�  +  ,9       .    ,  4� kH  ,� kH  ,� u  4� u  4� kH +  ,10      .    ,  4� (�  ,� (�  ,� kH  4� kH  4� (�      0    ,  % .�  L .�  L 6�  % 6�  % .�      0    ,  % F,  L F,  L M�  % M�  % F,      0    ,  % ]�  L ]�  L el  % el  % ]�      1    ,  ) *�  d *�  d iT  ) iT  ) *� +  ,11      +    ,  �� (�  p (�  p kH  �� kH  �� (�      *    ,  �( p     p     ��  �( ��  �( p +  ,13      ,    ,  �� !  � !  � s  �� s  �� !      +    ,  ,� (�  p (�  p kH  ,� kH  ,� (� +  ,12      +    ,  p  e�  ,�  e�  ,�  ��  p  ��  p  e� +  ,2       0    ,  L  kl  %  kl  %  s<  L  s<  L  kl      0    ,  L  ��  %  ��  %  ��  L  ��  L  ��      1    ,  d  g�  )  g�  )  ��  d  ��  d  g� +  ,1       .    ,  ,�  [�  4�  [�  4�  e�  ,�  e�  ,�  [� +  ,3       .    ,  ,�  ��  4�  ��  4�  �L  ,�  �L  ,�  �� +  ,4       .    ,  ,�  e�  4�  e�  4�  ��  ,�  ��  ,�  e�      .    ,  D\  [�  L,  [�  L,  e�  D\  e�  D\  [� +  ,5       .    ,  D\  ��  L,  ��  L,  �L  D\  �L  D\  �� +  ,6       .    ,  D\  e�  L,  e�  L,  ��  D\  ��  D\  e�      0    ,  S�  kl  [�  kl  [�  s<  S�  s<  S�  kl      0    ,  S�  ��  [�  ��  [�  ��  S�  ��  S�  ��      1    ,  P  g�  _�  g�  _�  ��  P  ��  P  g� +  ,7       .    ,  e�  s<  m`  s<  m`  }   e�  }   e�  s< +  ,8       .    ,  e�  ��  m`  ��  m`  �L  e�  �L  e�  �� +  ,9       .    ,  e�  }   m`  }   m`  ��  e�  ��  e�  }       0    ,  u0  ��  }   ��  }   ��  u0  ��  u0  ��      1    ,  qH  ~�  ��  ~�  ��  ��  qH  ��  qH  ~� +  ,10      +    <  a�  e�  a�  }   ��  }   ��  ��  p  ��  p  e�  a�  e�      )    <  y  N   y  e�  �L  e�  �L  ��      ��      N   y  N  +  ,12      -    <  ix  ]�  ix  u0  ��  u0  ��  �X  �  �X  �  ]�  ix  ]�      +    ,  m`  }   ��  }   ��  ��  m`  ��  m`  }  +  ,11   
  via    g�  ��   
  via    @  ��   
  via    Bh  ��   
  via    ��  ��      3    ,  ]�  ��  qH  ��  qH  �`  ]�  �`  ]�  ��      3    ,  |  ��  )  ��  )  �`  |  �`  |  ��      3    ,  8�  ��  L,  ��  L,  �`  8�  �`  8�  ��      3    ,  ��  ��  �p  ��  �p  �`  ��  �`  ��  ��      1    ,     ��  �( ��  �( ��     ��     ��      1    ,          �(      �(  '      '              0    ,  L,  |  S�  |  S�  L  L,  L  L,  |      0    ,  c�  |  kl  |  kl  L  c�  L  c�  |      0    ,  L, �t  S� �t  S� �D  L, �D  L, �t      0    ,  L �t  % �t  % �D  L �D  L �t      0    ,  {  |  ��  |  ��  L  {  L  {  |      0    ,  4�  |  <�  |  <�  L  4�  L  4�  |      0    ,  4� �t  <� �t  <� �D  4� �D  4� �t      0    ,  c� �t  kl �t  kl �D  c� �D  c� �t      0    ,  { �t  �� �t  �� �D  { �D  { �t      0    ,  L  |  %  |  %  L  L  L  L  |      0    ,  <� ��  D\ ��  D\ ��  <� ��  <� ��      0    ,  <� �4  D\ �4  D\ �  <� �  <� �4      0    ,  L  HD  %  HD  %  P  L  P  L  HD      0    ,  L  0�  %  0�  %  8�  L  8�  L  0�      0    ,  u0  _�  }   _�  }   g�  u0  g�  u0  _�      0    ,  u0  HD  }   HD  }   P  u0  P  u0  HD      0    ,  u0  0�  }   0�  }   8�  u0  8�  u0  0�   	   1      � $  ]� *�  ]� d  #( d  #( *�      1    ,  p  ��  '  ��  '  �l  p  �l  p  ��      1    ,  qH  '  ��  '  ��  kl  qH  kl  qH  '      1    ,  s<  kl  ��  kl  ��  ~�  s<  ~�  s<  kl   	   1      � 4  Y�  ��  Y�  ��  ��  ��  �� p  �� p  �� *�      1    ,  _�  ��  oT  ��  oT  �l  _�  �l  _�  ��      1    ,  :�  ��  J8  ��  J8  �l  :�  �l  :�  ��      1    ,  :� iT  FP iT  FP |�  :� |�  :� iT      1    ,  8� |�  HD |�  HD ��  8� ��  8� |�      1    ,  d  S�  '  S�  '  g�  d  g�  d  S�      1    ,  d  '  )  '  )  S�  d  S�  d  '      +    ,  p ��  �� ��  �� �   p �   p ��      +    ,  p  �  ��  �  ��  #(  p  #(  p  �      +    ,  6� z�  J8 z�  J8 ��  6� ��  6� z�      +    ,  8� kH  HD kH  HD z�  8� z�  8� kH      +    ,  p  U�  )  U�  )  e�  p  e�  p  U�      +    ,  p  #(  *�  #(  *�  U�  p  U�  p  #(      +    ,  qH  m`  ��  m`  ��  }   qH  }   qH  m`      +    ,  oT  #(  ��  #(  ��  m`  oT  m`  oT  #(      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      ,    ,  �  *�  2�  *�  2�  ]�  �  ]�  �  *�      ,    <  g�  *�  ��  *�  ��  u0  ix  u0  ix  ]�  g�  ]�  g�  *�      -    ,  � ��  �� ��  �� ��  � ��  � ��      -    ,  .� s  R s  R ��  .� ��  .� s      )    ,          �(      �(  ��      ��              *    ,     p  �( p  �( ��     ��     p      .    ,  8�  ��  L,  ��  L,  �`  8�  �`  8�  ��   	   .      � $  P   P �  HD �  HD  �L   	   .      �   oT   oT  �L  e�  �L   	   .      � $  0�   0� �  % �  %  �`      .    ,  ]�  ��  qH  ��  qH  �`  ]�  �`  ]�  ��      .    ,  |  ��  )  ��  )  �`  |  �`  |  ��   	   .      �   %  ��  %  �L  4�  �L      /    ,  c�  ܴ  kl  ܴ  kl  �  c�  �  c�  ܴ      /    ,  >�  ܴ  FP  ܴ  FP  �  >�  �  >�  ܴ      /    ,  X  ܴ  #(  ܴ  #(  �  X  �  X  ܴ              P  � GND  +  ,1               P �8 VDD  +  ,1               @  �� A1 +  ,1               Bh  �� A0 +  ,1               g�  �� B0 +  ,1               ��  �� Y  +  ,1       �    ,          �(      �( ��     ��                      P  � GND               P �8 VDD               @  �� A1              Bh  �� A0              g�  �� B0              ��  �� Y      �     $� 	   /  
aoi221    0    ,  �� #  { #  { *�  �� *�  �� #      0    ,  �� :t  { :t  { BD  �� BD  �� :t      0    ,  �� Q�  { Q�  { Y�  �� Y�  �� Q�      0    ,  �� iT  { iT  { q$  �� q$  �� iT      1    ,  ��   w$   w$ u  �� u  ��  +  ,1       .    ,  s< d  kl d  kl (  s< (  s< d +  ,3       .    ,  s< w   kl w   kl ��  s< ��  s< w  +  ,4       .    ,  s< (  kl (  kl w   s< w   s< (      0    ,  c� #  [� #  [� *�  c� *�  c� #      0    ,  c� :t  [� :t  [� BD  c� BD  c� :t      0    ,  c� Q�  [� Q�  [� Y�  c� Y�  c� Q�      0    ,  c� iT  [� iT  [� q$  c� q$  c� iT      1    ,  g�   W�   W� u  g� u  g�  +  ,5       .    ,  S� d  L, d  L, (  S� (  S� d +  ,6       .    ,  S� w   L, w   L, ��  S� ��  S� w  +  ,7       .    ,  S� (  L, (  L, w   S� w   S� (      0    ,  D\ #  <� #  <� *�  D\ *�  D\ #      0    ,  D\ :t  <� :t  <� BD  D\ BD  D\ :t      0    ,  D\ Q�  <� Q�  <� Y�  D\ Y�  D\ Q�      0    ,  D\ iT  <� iT  <� q$  D\ q$  D\ iT      1    ,  HD   8�   8� u  HD u  HD  +  ,8       .    ,  4� d  ,� d  ,� (  4� (  4� d +  ,9       .    ,  4� w   ,� w   ,� ��  4� ��  4� w  +  ,10      .    ,  4� (  ,� (  ,� w   4� w   4� (      0    ,  % #  L #  L *�  % *�  % #      0    ,  % :t  L :t  L BD  % BD  % :t      0    ,  % Q�  L Q�  L Y�  % Y�  % Q�      0    ,  % iT  L iT  L q$  % q$  % iT      1    ,  )   d   d u  ) u  )  +  ,11      +    ,  �� (  p (  p w   �� w   �� (      *    ,  �( �     �     �p  �( �p  �( � +  ,13      ,    ,  �� X  � X  � ~�  �� ~�  �� X      +    ,  �� (  s< (  s< w   �� w   �� ( +  ,2       +    ,  ,� (  p (  p w   ,� w   ,� ( +  ,12      +    ,  �p (  �� (  �� w   �p w   �p ( +  ,2       0    ,  �L #  � #  � *�  �L *�  �L #      0    ,  �L :t  � :t  � BD  �L BD  �L :t      0    ,  �L Q�  � Q�  � Y�  �L Y�  �L Q�      0    ,  �L iT  � iT  � q$  �L q$  �L iT      1    ,  �d   �   � u  �d u  �d  +  ,1       .    ,  �� d  �� d  �� (  �� (  �� d +  ,3       .    ,  �� w   �� w   �� ��  �� ��  �� w  +  ,4       .    ,  �� (  �� (  �� w   �� w   �� (      0    ,  �� #  �\ #  �\ *�  �� *�  �� #      0    ,  �� :t  �\ :t  �\ BD  �� BD  �� :t      0    ,  �� Q�  �\ Q�  �\ Y�  �� Y�  �� Q�      0    ,  �� iT  �\ iT  �\ q$  �� q$  �� iT      1    ,  ��   �D   �D u  �� u  ��  +  ,5       .    ,  �, d  �� d  �� (  �, (  �, d +  ,6       .    ,  �, w   �� w   �� ��  �, ��  �, w  +  ,7       .    ,  �, (  �� (  �� w   �, w   �, (      0    ,  �� #  �� #  �� *�  �� *�  �� #      0    ,  �� :t  �� :t  �� BD  �� BD  �� :t      0    ,  �� Q�  �� Q�  �� Y�  �� Y�  �� Q�      0    ,  �� iT  �� iT  �� q$  �� q$  �� iT      1    ,  ��   �   � u  �� u  ��  +  ,8       +    ,  �p (  �x (  �x w   �p w   �p (      *    ,  }  �  �� �  �� �p  }  �p  }  � +  ,10      ,    ,  �� X  �H X  �H ~�  �� ~�  �� X      +    ,  �� (  �x (  �x w   �� w   �� ( +  ,9       +    ,  p  }   ,�  }   ,�  ��  p  ��  p  }  +  ,2       0    ,  L  ��  %  ��  %  ��  L  ��  L  ��      1    ,  d  ~�  )  ~�  )  ��  d  ��  d  ~� +  ,1       .    ,  ,�  s<  4�  s<  4�  }   ,�  }   ,�  s< +  ,3       .    ,  ,�  ��  4�  ��  4�  �L  ,�  �L  ,�  �� +  ,4       .    ,  ,�  }   4�  }   4�  ��  ,�  ��  ,�  }       0    ,  >�  kl  FP  kl  FP  s<  >�  s<  >�  kl      0    ,  >�  ��  FP  ��  FP  ��  >�  ��  >�  ��      1    ,  :�  g�  J8  g�  J8  ��  :�  ��  :�  g� +  ,5       .    ,  N   [�  U�  [�  U�  e�  N   e�  N   [� +  ,6       .    ,  N   ��  U�  ��  U�  �L  N   �L  N   �� +  ,7       .    ,  N   e�  U�  e�  U�  ��  N   ��  N   e�      .    ,  e�  [�  m`  [�  m`  e�  e�  e�  e�  [� +  ,8       .    ,  e�  ��  m`  ��  m`  �L  e�  �L  e�  �� +  ,9       .    ,  e�  e�  m`  e�  m`  ��  e�  ��  e�  e�      0    ,  w$  c�  ~�  c�  ~�  kl  w$  kl  w$  c�      0    ,  w$  {  ~�  {  ~�  ��  w$  ��  w$  {      1    ,  s<  _�  ��  _�  ��  ��  s<  ��  s<  _� +  ,10      .    ,  ��  S�  ��  S�  ��  ]�  ��  ]�  ��  S� +  ,11      .    ,  ��  ��  ��  ��  ��  �L  ��  �L  ��  �� +  ,12      .    ,  ��  ]�  ��  ]�  ��  ��  ��  ��  ��  ]�      .    ,  �4  S�  �  S�  �  ]�  �4  ]�  �4  S� +  ,13      .    ,  �4  ��  �  ��  �  �L  �4  �L  �4  �� +  ,14      .    ,  �4  ]�  �  ]�  �  ��  �4  ��  �4  ]�      0    ,  ��  kl  ��  kl  ��  s<  ��  s<  ��  kl      0    ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��      1    ,  ��  g�  ��  g�  ��  ��  ��  ��  ��  g� +  ,15      +    \  ��  ]�  ��  e�  ��  e�  ��  ��  p  ��  p  }   8�  }   8�  e�  qH  e�  qH  ]�  ��  ]�      )    \  �  FP  �  N   ��  N   ��  ��      ��      e�  !4  e�  !4  N   Y�  N   Y�  FP  �  FP +  ,17      -    \  �t  U�  �t  ]�  �P  ]�  �P  �X  �  �X  �  u0  0�  u0  0�  ]�  ix  ]�  ix  U�  �t  U�      +    <  ��  ]�  ��  e�  ��  e�  ��  ��  �  ��  �  ]�  ��  ]� +  ,16   
  via  �  B�         HD  �   
  via  �  B�         ��  �   
  via  �  B�         ��  �   
  via  �  B�         ��  �   
  via  �  B�         kl  �   
  via  �  B�         %  �      1    ,     ��  �� ��  �� ��     ��     ��      1    ,          ��      ��  '      '              1    ,     ��  �� ��  �� ��     ��     ��      1    ,          ��      ��  '      '              3    ,  �   �P  ި  �P  ި  ��  �   ��  �   �P      3    ,  >�  �P  R  �P  R  ��  >�  ��  >�  �P      3    ,  a�  �P  u0  �P  u0  ��  a�  ��  a�  �P      3    ,  ��  �P  ��  �P  ��  ��  ��  ��  ��  �P      3    ,  ��  �P  �X  �P  �X  ��  ��  ��  ��  �P      3    ,  X  �P  .�  �P  .�  ��  X  ��  X  �P      /    ,  ��  �,  ��  �,  ��  ��  ��  ��  ��  �,      /    ,  ��  �,  ��  �,  ��  ��  ��  ��  ��  �,      /    ,  g�  �,  oT  �,  oT  ��  g�  ��  g�  �,      /    ,  FP  �,  N   �,  N   ��  FP  ��  FP  �,      /    ,  #(  �,  *�  �,  *�  ��  #(  ��  #(  �,   	   .      � $  ��  �L  ��  ��  ��  ��  �� d      .    ,  L  �P  0�  �P  0�  ��  L  ��  L  �P   	   .      �   0� d  0�  �L   	   .      �   P d  P  �L  U�  �L   	   .      �   e�  �L  oT  �L  oT d      .    ,  �   �P  ި  �P  ި  ��  �   ��  �   �P      .    ,  ��  �P  ��  �P  ��  ��  ��  ��  ��  �P      .    ,  a�  �P  u0  �P  u0  ��  a�  ��  a�  �P      .    ,  @t  �P  S�  �P  S�  ��  @t  ��  @t  �P   	   .      �   � d  �  �L  �4  �L      *    ,     �  �� �  �� ��     ��     �      )    ,          ��      ��  ��      ��              ,    ,  �  �  �H  �  �H  *�  �  *�  �  �      ,    <  �  *�  2�  *�  2�  ]�  0�  ]�  0�  u0  �  u0  �  *�      ,    ,  ix  *�  ��  *�  ��  U�  ix  U�  ix  *�      -    ,  � ��  �H ��  �H ��  � ��  � ��      -    ,  �� ~�  � ~�  � ��  �� ��  �� ~�      +    ,  p  �  �x  �  �x  #(  p  #(  p  �      +    ,  p ��  �x ��  �x �   p �   p ��      +    ,  p  m`  )  m`  )  }   p  }   p  m`      +    ,  p  #(  *�  #(  *�  m`  p  m`  p  #(      +    ,  qH  N   ��  N   ��  ]�  qH  ]�  qH  N       +    ,  qH  #(  ��  #(  ��  N   qH  N   qH  #(      +    ,  �� ��  �8 ��  �8 ��  �� ��  �� ��      +    ,  �� w   �D w   �D ��  �� ��  �� w    	   1      � $  }  u  }  �p  Bh �p  Bh u      1    ,  @  �D  .�  �D  .�  ��  @  ��  @  �D   	   1      � $  #(   #(  �<  ��  �<  ��  ��   	   1      �   ��  �P  ��  ��   	   1      � $  �@   �@ �  a� �  a�    	   1      � $  �(   �( �  �� �  ��    	   1      � $  D\  ��  D\  ��  ��  ��  ��  ��      1    ,  �  �D  ܴ  �D  ܴ  ��  �  ��  �  �D      1    ,  ��  �D  ��  �D  ��  ��  ��  ��  ��  �D      1    ,  c�  �D  s<  �D  s<  ��  c�  ��  c�  �D      1    ,  Bh  �D  R  �D  R  ��  Bh  ��  Bh  �D      1    ,  d  '  )  '  )  kl  d  kl  d  '      1    ,  d  kl  '  kl  '  ~�  d  ~�  d  kl      1    ,  s<  L,  ��  L,  ��  _�  s<  _�  s<  L,      1    ,  s<  '  ��  '  ��  L,  s<  L,  s<  '      1    ,  �� u  �P u  �P ��  �� ��  �� u      1    ,  �� ��  �D ��  �D ��  �� ��  �� ��      0    ,  {  |  ��  |  ��  L  {  L  {  |      0    ,  c�  |  kl  |  kl  L  c�  L  c�  |      0    ,  �|  |  �L  |  �L  L  �|  L  �|  |      0    ,  L,  |  S�  |  S�  L  L,  L  L,  |      0    ,  L, �t  S� �t  S� �D  L, �D  L, �t      0    ,  c� �t  kl �t  kl �D  c� �D  c� �t      0    ,  ��  |  ��  |  ��  L  ��  L  ��  |      0    ,  �\  |  �,  |  �,  L  �\  L  �\  |      0    ,  ��  |  ��  |  ��  L  ��  L  ��  |      0    ,  4�  |  <�  |  <�  L  4�  L  4�  |      0    ,  4� �t  <� �t  <� �D  4� �D  4� �t      0    ,  L  |  %  |  %  L  L  L  L  |      0    ,  �� �t  �� �t  �� �D  �� �D  �� �t      0    ,  �\ �t  �, �t  �, �D  �\ �D  �\ �t      0    ,  �� �t  �� �t  �� �D  �� �D  �� �t      0    ,  �| �t  �L �t  �L �D  �| �D  �| �t      0    ,  { �t  �� �t  �� �D  { �D  { �t      0    ,  L �t  % �t  % �D  L �D  L �t      0    ,  L  _�  %  _�  %  g�  L  g�  L  _�      0    ,  L  HD  %  HD  %  P  L  P  L  HD      0    ,  L  0�  %  0�  %  8�  L  8�  L  0�      0    ,  w$  @t  ~�  @t  ~�  HD  w$  HD  w$  @t      0    ,  �� �|  �\ �|  �\ �L  �� �L  �� �|              ~�  � GND  +  ,1               ~� �8 VDD  +  ,1               ��  � A1 +  ,1               ��  � A0 +  ,1               %  � C0 +  ,1               kl  � B1 +  ,1               HD  � B0 +  ,1               ��  � Y  +  ,1       �    ,          ��      �� ��     ��                      ~�  � GND               ~� �8 VDD               ��  � A1              ��  � A0              %  � C0              kl  � B1              HD  � B0              ��  � Y      �   
 ' � 	   /  ao22    0    ,  L   %   % &�  L &�  L       0    ,  L 6�  % 6�  % >\  L >\  L 6�      0    ,  L M�  % M�  % U�  L U�  L M�      1    ,  d 4  ) 4  ) Y�  d Y�  d 4 +  ,1       .    ,  ,� |  4� |  4� @  ,� @  ,� | +  ,3       .    ,  ,� [�  4� [�  4� el  ,� el  ,� [� +  ,4       .    ,  ,� @  4� @  4� [�  ,� [�  ,� @      0    ,  <�   D\   D\ &�  <� &�  <�       0    ,  <� 6�  D\ 6�  D\ >\  <� >\  <� 6�      0    ,  <� M�  D\ M�  D\ U�  <� U�  <� M�      1    ,  8� 4  HD 4  HD Y�  8� Y�  8� 4 +  ,5       .    ,  L, |  S� |  S� @  L, @  L, | +  ,6       .    ,  L, [�  S� [�  S� el  L, el  L, [� +  ,7       .    ,  L, @  S� @  S� [�  L, [�  L, @      0    ,  [�   c�   c� &�  [� &�  [�       0    ,  [� 6�  c� 6�  c� >\  [� >\  [� 6�      0    ,  [� M�  c� M�  c� U�  [� U�  [� M�      1    ,  W� 4  g� 4  g� Y�  W� Y�  W� 4 +  ,8       .    ,  kl |  s< |  s< @  kl @  kl | +  ,9       .    ,  kl [�  s< [�  s< el  kl el  kl [� +  ,10      .    ,  kl @  s< @  s< [�  kl [�  kl @      0    ,  {   ��   �� &�  { &�  {       0    ,  { 6�  �� 6�  �� >\  { >\  { 6�      0    ,  { M�  �� M�  �� U�  { U�  { M�      1    ,  w$ 4  �� 4  �� Y�  w$ Y�  w$ 4 +  ,11      .    ,  �� |  �| |  �| @  �� @  �� | +  ,12      .    ,  �� [�  �| [�  �| el  �� el  �� [� +  ,13      .    ,  �� @  �| @  �| [�  �� [�  �� @      0    ,  �L   �   � &�  �L &�  �L       0    ,  �L 6�  � 6�  � >\  �L >\  �L 6�      0    ,  �L M�  � M�  � U�  �L U�  �L M�      1    ,  �d 4  � 4  � Y�  �d Y�  �d 4 +  ,14      .    ,  �� |  �� |  �� @  �� @  �� | +  ,15      .    ,  �� D8  �� D8  �� M�  �� M�  �� D8 +  ,16      .    ,  �� @  �� @  �� D8  �� D8  �� @      0    ,  ��   �P   �P &�  �� &�  ��       0    ,  �� 6�  �P 6�  �P >\  �� >\  �� 6�      1    ,  �� 4  �8 4  �8 BD  �� BD  �� 4 +  ,17      +    <  �, @  �, D8  �� D8  �� [�  p [�  p @  �, @      *    <  �� �  �� [�  �h [�  �h s     s     �  �� � +  ,19      ,    <  �� p  �� L  �� L  �� cx  � cx  � p  �� p      +    ,  p @  ,� @  ,� [�  p [�  p @ +  ,2       +    ,  �� @  �, @  �, D8  �� D8  �� @ +  ,18      +    ,  @  e�  4�  e�  4�  ��  @  ��  @  e� +  ,2       0    ,  %  kl  ,�  kl  ,�  s<  %  s<  %  kl      0    ,  %  ��  ,�  ��  ,�  ��  %  ��  %  ��      1    ,  !4  g�  0�  g�  0�  ��  !4  ��  !4  g� +  ,1       .    ,  4�  [�  <�  [�  <�  e�  4�  e�  4�  [� +  ,3       .    ,  4�  ��  <�  ��  <�  �L  4�  �L  4�  �� +  ,4       .    ,  4�  e�  <�  e�  <�  ��  4�  ��  4�  e�      .    ,  L,  [�  S�  [�  S�  e�  L,  e�  L,  [� +  ,5       .    ,  L,  ��  S�  ��  S�  �L  L,  �L  L,  �� +  ,6       .    ,  L,  e�  S�  e�  S�  ��  L,  ��  L,  e�      0    ,  [�  kl  c�  kl  c�  s<  [�  s<  [�  kl      0    ,  [�  ��  c�  ��  c�  ��  [�  ��  [�  ��      1    ,  W�  g�  g�  g�  g�  ��  W�  ��  W�  g� +  ,7       .    ,  kl  [�  s<  [�  s<  e�  kl  e�  kl  [� +  ,8       .    ,  kl  ��  s<  ��  s<  �L  kl  �L  kl  �� +  ,9       .    ,  kl  e�  s<  e�  s<  ��  kl  ��  kl  e�      .    ,  ��  [�  ��  [�  ��  e�  ��  e�  ��  [� +  ,10      .    ,  ��  ��  ��  ��  ��  �L  ��  �L  ��  �� +  ,11      .    ,  ��  e�  ��  e�  ��  ��  ��  ��  ��  e�      0    ,  �|  kl  �L  kl  �L  s<  �|  s<  �|  kl      0    ,  �|  ��  �L  ��  �L  ��  �|  ��  �|  ��      1    ,  ��  g�  �4  g�  �4  ��  ��  ��  ��  g� +  ,12      .    ,  �  s<  ��  s<  ��  }   �  }   �  s< +  ,13      .    ,  �  ��  ��  ��  ��  �L  �  �L  �  �� +  ,14      .    ,  �  }   ��  }   ��  ��  �  ��  �  }       0    ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��      1    ,  ��  ~�  �h  ~�  �h  ��  ��  ��  ��  ~� +  ,15      +    <  �(  e�  �(  }   �\  }   �\  ��  @  ��  @  e�  �(  e�      )    <  ��  N   ��  e�  ��  e�  ��  ��  �  ��  �  N   ��  N  +  ,17      -    <  ��  ]�  ��  u0  �,  u0  �,  �X  p  �X  p  ]�  ��  ]�      +    ,  ��  }   �\  }   �\  ��  ��  ��  ��  }  +  ,16   
  via    p  �   
  via    ��  �   
  via    �8  �   
  via    :�  �   
  via    ]�  �      1    ,     ��  �� ��  �� ��     ��     ��      1    ,          ��      ��  '      '              1    ,     ��  �� ��  �� ��     ��     ��      1    ,          ��      ��  '      '              3    ,  �t  �P  ��  �P  ��  ��  �t  ��  �t  �P      3    ,  {  �P  ��  �P  ��  ��  {  ��  {  �P      3    ,  0�  �P  D\  �P  D\  ��  0�  ��  0�  �P      3    ,  �  �P  !4  �P  !4  ��  �  ��  �  �P      3    ,  S�  �P  g�  �P  g�  ��  S�  ��  S�  �P      /    ,  6�  �,  >�  �,  >�  ��  6�  ��  6�  �,      /    ,  ��  �T  �p  �T  �p  �$  ��  �$  ��  �T      /    ,  ��  �,  ��  �,  ��  ��  ��  ��  ��  �,      /    ,  �  �,  X  �,  X  ��  �  ��  �  �,      /    ,  Y�  �,  a�  �,  a�  ��  Y�  ��  Y�  �,      /    ,  �  �,  ��  �,  ��  ��  �  ��  �  �,   	   .      � $  P |  P  �   W�  �   W�  ��   	   .      �   �� |  ��  ��      .    ,  {  �P  ��  �P  ��  ��  {  ��  {  �P   	   .      � $  oT |  oT  �   w$  �   w$  �      .    ,  S�  �P  g�  �P  g�  ��  S�  ��  S�  �P   	   .      � $  oT  �L  oT  ��  c�  ��  c�  �P      .    ,  �  �P  !4  �P  !4  ��  �  ��  �  �P   	   .      �   ��  �L  ��  �P      .    ,  0�  �P  D\  �P  D\  ��  0�  ��  0�  �P      .    ,  ��  �x  �L  �x  �L  �   ��  �   ��  �x   	   .      �   <�  �L  L  �L  L  �P   	   .      � $  P  �L  P  ��  @t  ��  @t  �P   	   .      �   �� |  ��  �    	   .      �   L  ��  L |  4� |      .    ,  �(  �P  ��  �P  ��  ��  �(  ��  �(  �P   	   .      �   ��  �P  ��  �L  �  �L      *    ,     �  �� �  �� ��     ��     �      )    ,          ��      ��  ��      ��              -    ,  � ��  �� ��  �� ��  � ��  � ��      -    ,  �� cx  �� cx  �� ��  �� ��  �� cx      -    ,  � cx  2� cx  2� ��  � ��  � cx      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      ,    ,  ��  *�  ��  *�  ��  ]�  ��  ]�  ��  *�      ,    ,  p  *�  :�  *�  :�  ]�  p  ]�  p  *�      0    ,  �  |  ��  |  ��  L  �  L  �  |      0    ,  d  |  !4  |  !4  L  d  L  d  |      0    ,  0�  |  8�  |  8�  L  0�  L  0�  |      0    ,  HD  |  P  |  P  L  HD  L  HD  |      0    ,  _�  |  g�  |  g�  L  _�  L  _�  |      0    ,  w$  |  ~�  |  ~�  L  w$  L  w$  |      0    ,  ��  |  �d  |  �d  L  ��  L  ��  |      0    ,  �t  |  �D  |  �D  L  �t  L  �t  |      0    ,  �t �t  �D �t  �D �D  �t �D  �t �t      0    ,  � �t  �� �t  �� �D  � �D  � �t      0    ,  �� �t  �d �t  �d �D  �� �D  �� �t      0    ,  w$ �t  ~� �t  ~� �D  w$ �D  w$ �t      0    ,  _� �t  g� �t  g� �D  _� �D  _� �t      0    ,  HD �t  P �t  P �D  HD �D  HD �t      0    ,  0� �t  8� �t  8� �D  0� �D  0� �t      0    ,  d �t  !4 �t  !4 �D  d �D  d �t      0    ,  �L q$  � q$  � x�  �L x�  �L q$      0    ,  �L ��  � ��  � �d  �L �d  �L ��      0    ,  �L �  � �  � ��  �L ��  �L �      0    ,  L q$  % q$  % x�  L x�  L q$      0    ,  L ��  % ��  % �d  L �d  L ��      0    ,  L �  % �  % ��  L ��  L �      0    ,  �|  HD  �L  HD  �L  P  �|  P  �|  HD      0    ,  �|  0�  �L  0�  �L  8�  �|  8�  �|  0�      0    ,  %  HD  ,�  HD  ,�  P  %  P  %  HD      0    ,  %  0�  ,�  0�  ,�  8�  %  8�  %  0�      +    ,  �  �  �   �  �   #(  �  #(  �  �      +    ,  � ��  �  ��  �  �   � �   � ��      +    ,  �p kH  �� kH  �� ��  �p ��  �p kH      +    ,  �d [�  �� [�  �� kH  �d kH  �d [�      +    ,  p kH  *� kH  *� ��  p ��  p kH      +    ,  p [�  ) [�  ) kH  p kH  p [�      +    ,  ��  U�  �(  U�  �(  e�  ��  e�  ��  U�      +    ,  ��  #(  �(  #(  �(  U�  ��  U�  ��  #(      +    ,  @  #(  2�  #(  2�  U�  @  U�  @  #(      +    ,  @  U�  0�  U�  0�  e�  @  e�  @  U�      1    ,  �  �D  ��  �D  ��  ��  �  ��  �  �D   	   1      � $  �(  ��  �(  ��  a�  ��  a�  ��      1    ,  2�  �D  Bh  �D  Bh  ��  2�  ��  2�  �D   	   1      � $  }  Y�  }  s  Bh s  Bh Y�   	   1      �   �P &�  �P  ��   	   1      � $  a� 4  a� 	�  �� 	�  ��  ��      1    ,  �  �D  @  �D  @  ��  �  ��  �  �D   	   1      �   ��  �H  <�  �H  <�  ��      1    ,  ��  �l  �X  �l  �X  �  ��  �  ��  �l      1    ,  U�  �D  e�  �D  e�  ��  U�  ��  U�  �D      1    ,  }   �D  ��  �D  ��  ��  }   ��  }   �D      1    ,  �X Y�  � Y�  � m<  �X m<  �X Y�      1    ,  �d m<  � m<  � ��  �d ��  �d m<      1    ,  d m<  ) m<  ) ��  d ��  d m<      1    ,  d Y�  ' Y�  ' m<  d m<  d Y�      1    ,  ��  S�  �4  S�  �4  g�  ��  g�  ��  S�      1    ,  ��  '  �4  '  �4  S�  ��  S�  ��  '      1    ,  !4  '  0�  '  0�  S�  !4  S�  !4  '      1    ,  !4  S�  .�  S�  .�  g�  !4  g�  !4  S�              pN  � GND  +  ,1               pN �8 VDD  +  ,1               p  � A1 +  ,1               �8  � Y  +  ,1               ��  � B1 +  ,1               :�  � A0 +  ,1               ]�  � B0 +  ,1       �    ,          ��      �� ��     ��                      p  � A1              pN  � GND               pN �8 VDD               �8  � Y               ��  � B1              :�  � A0              ]�  � B0     �    ' %� 	   0 : 
oai22     0    ,  % �  ,� �  ,� |  % |  % �      0    ,  %   ,�   ,� &�  % &�  %       0    ,  % 6�  ,� 6�  ,� >\  % >\  % 6�      0    ,  % M�  ,� M�  ,� U�  % U�  % M�      0    ,  % el  ,� el  ,� m<  % m<  % el      1    ,  !4 �  0� �  0� q$  !4 q$  !4 � +  ,1       .    ,  4�  �  <�  �  <� �  4� �  4�  � +  ,3       .    ,  4� s  <� s  <� |�  4� |�  4� s +  ,4       .    ,  4� �  <� �  <� s  4� s  4� �      .    ,  L,  �  S�  �  S� �  L, �  L,  � +  ,5       .    ,  L, s  S� s  S� |�  L, |�  L, s +  ,6       .    ,  L, �  S� �  S� s  L, s  L, �      0    ,  [� �  c� �  c� |  [� |  [� �      0    ,  [�   c�   c� &�  [� &�  [�       0    ,  [� 6�  c� 6�  c� >\  [� >\  [� 6�      0    ,  [� M�  c� M�  c� U�  [� U�  [� M�      0    ,  [� el  c� el  c� m<  [� m<  [� el      1    ,  W� �  g� �  g� q$  W� q$  W� � +  ,7       .    ,  kl  �  s<  �  s< �  kl �  kl  � +  ,8       .    ,  kl s  s< s  s< |�  kl |�  kl s +  ,9       .    ,  kl �  s< �  s< s  kl s  kl �      .    ,  ��  �  ��  �  �� �  �� �  ��  � +  ,10      .    ,  �� s  �� s  �� |�  �� |�  �� s +  ,11      .    ,  �� �  �� �  �� s  �� s  �� �      0    ,  �| �  �L �  �L |  �| |  �| �      0    ,  �|   �L   �L &�  �| &�  �|       0    ,  �| 6�  �L 6�  �L >\  �| >\  �| 6�      0    ,  �| M�  �L M�  �L U�  �| U�  �| M�      0    ,  �| el  �L el  �L m<  �| m<  �| el      1    ,  �� �  �4 �  �4 q$  �� q$  �� � +  ,12      +    ,  @ �  �( �  �( s  @ s  @ �      *    ,  �  �`  ��  �`  �� ��  � ��  �  �` +  ,14      ,    ,  p  �   ��  �   �� z�  p z�  p  �       +    ,  @ �  4� �  4� s  @ s  @ � +  ,2       +    ,  �� �  �( �  �( s  �� s  �� � +  ,13      0    ,  �  ]�  �L  ]�  �L  e�  �  e�  �  ]�      0    ,  �  u0  �L  u0  �L  }   �  }   �  u0      1    ,  �  Y�  �d  Y�  �d  ��  �  ��  �  Y� +  ,1       .    ,  �|  N   ��  N   ��  W�  �|  W�  �|  N  +  ,3       .    ,  �|  ��  ��  ��  ��  ��  �|  ��  �|  �� +  ,4       .    ,  �|  W�  ��  W�  ��  ��  �|  ��  �|  W�      0    ,  ��  ]�  {  ]�  {  e�  ��  e�  ��  ]�      0    ,  ��  u0  {  u0  {  }   ��  }   ��  u0      1    ,  ��  Y�  w$  Y�  w$  ��  ��  ��  ��  Y� +  ,5       .    ,  s<  N   kl  N   kl  W�  s<  W�  s<  N  +  ,6       .    ,  s<  ��  kl  ��  kl  ��  s<  ��  s<  �� +  ,7       .    ,  s<  W�  kl  W�  kl  ��  s<  ��  s<  W�      0    ,  c�  ]�  [�  ]�  [�  e�  c�  e�  c�  ]�      0    ,  c�  u0  [�  u0  [�  }   c�  }   c�  u0      1    ,  g�  Y�  W�  Y�  W�  ��  g�  ��  g�  Y� +  ,8       .    ,  S�  N   L,  N   L,  W�  S�  W�  S�  N  +  ,9       .    ,  S�  ��  L,  ��  L,  ��  S�  ��  S�  �� +  ,10      .    ,  S�  W�  L,  W�  L,  ��  S�  ��  S�  W�      0    ,  D\  ]�  <�  ]�  <�  e�  D\  e�  D\  ]�      0    ,  D\  u0  <�  u0  <�  }   D\  }   D\  u0      1    ,  HD  Y�  8�  Y�  8�  ��  HD  ��  HD  Y� +  ,11      .    ,  4�  N   ,�  N   ,�  W�  4�  W�  4�  N  +  ,12      .    ,  4�  ��  ,�  ��  ,�  ��  4�  ��  4�  �� +  ,13      .    ,  4�  W�  ,�  W�  ,�  ��  4�  ��  4�  W�      0    ,  %  ]�  L  ]�  L  e�  %  e�  %  ]�      0    ,  %  u0  L  u0  L  }   %  }   %  u0      1    ,  )  Y�  d  Y�  d  ��  )  ��  )  Y� +  ,14      +    ,  ��  W�  p  W�  p  ��  ��  ��  ��  W�      )    ,  �h  @t      @t      �L  �h  �L  �h  @t +  ,16      -    ,  ��  P  �  P  �  ��  ��  ��  ��  P      +    ,  ,�  W�  p  W�  p  ��  ,�  ��  ,�  W� +  ,15      +    ,  ��  W�  �|  W�  �|  ��  ��  ��  ��  W� +  ,2    
  via    d  �   
  via    ��  �   
  via    <�  �   
  via    _�  �   
  via    �  �      3    ,  U�  �P  ix  �P  ix  ��  U�  ��  U�  �P      3    ,  y  �P  ��  �P  ��  ��  y  ��  y  �P      3    ,  �  �P  #(  �P  #(  ��  �  ��  �  �P      3    ,  2�  �P  FP  �P  FP  ��  2�  ��  2�  �P      3    ,  �@  �P  ��  �P  ��  ��  �@  ��  �@  �P      1    ,          �h      �h  '      '              1    ,     ��  �h ��  �h ��     ��     ��      �    ,          �h      �h ��     ��              .    ,  2�  �P  FP  �P  FP  ��  2�  ��  2�  �P      .    ,  �@  �P  ��  �P  ��  ��  �@  ��  �@  �P      .    ,  y  �P  ��  �P  ��  ��  y  ��  y  �P      .    ,  �  �P  #(  �P  #(  ��  �  ��  �  �P   	   .      �   ��  �$  �(  �$  �(  ��   	   .      � $  }   ��  }   ��  oT  ��  oT  �   	   .      �   <�  �$  @  �$  @  ��   	   .      � $  Bh  ��  Bh  ��  P  ��  P  �   	   .      � $  Bh  �P  Bh  �  P  �  P  ��   	   .      � $  oT  ��  oT  ��  }   ��  }   �P   	   .      �   4�  ��  @  ��  @  �P   	   .      � $  �(  �P  �(  ��  ��  ��  ��  ��      /    ,  �  �,  ��  �,  ��  ��  �  ��  �  �,      /    ,  ~�  �,  ��  �,  ��  ��  ~�  ��  ~�  �,      /    ,  8�  �,  @t  �,  @t  ��  8�  ��  8�  �,      /    ,  |  �,  L  �,  L  ��  |  ��  |  �,      )    ,          �h      �h  ��      ��              *    ,      �`  �h  �`  �h ��     ��      �`      -    ,  � ��  �� ��  �� ��  � ��  � ��      -    ,  p z�  :� z�  :� ��  p ��  p z�      -    ,  �� z�  �� z�  �� ��  �� ��  �� z�      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      ,    ,  m`  *�  ��  *�  ��  P  m`  P  m`  *�      0    ,  | �t  L �t  L �D  | �D  | �t      0    ,  ,� �t  4� �t  4� �D  ,� �D  ,� �t      0    ,  D\ �t  L, �t  L, �D  D\ �D  D\ �t      0    ,  [� �t  c� �t  c� �D  [� �D  [� �t      0    ,  s< �t  { �t  { �D  s< �D  s< �t      0    ,  �� �t  �| �t  �| �D  �� �D  �� �t      0    ,  � �t  �� �t  �� �D  � �D  � �t      0    ,  �  |  ��  |  ��  L  �  L  �  |      0    ,  ��  |  �|  |  �|  L  ��  L  ��  |      0    ,  s<  |  {  |  {  L  s<  L  s<  |      0    ,  [�  |  c�  |  c�  L  [�  L  [�  |      0    ,  D\  |  L,  |  L,  L  D\  L  D\  |      0    ,  ,�  |  4�  |  4�  L  ,�  L  ,�  |      0    ,  |  |  L  |  L  L  |  L  |  |      0    ,  % �  ,� �  ,� ��  % ��  % �      0    ,  % ��  ,� ��  ,� �p  % �p  % ��      0    ,  �| �  �L �  �L ��  �| ��  �| �      0    ,  �| ��  �L ��  �L �p  �| �p  �| ��      0    ,  {  :�  ��  :�  ��  Bh  {  Bh  {  :�      1    ,  4�  �D  D\  �D  D\  ��  4�  ��  4�  �D      1    ,  �4  �D  ��  �D  ��  ��  �4  ��  �4  �D      1    ,  {  �D  ��  �D  ��  ��  {  ��  {  �D      1    ,  �  �D  !4  �D  !4  ��  �  ��  �  �D   	   1      � $  _�  �P  _�  ��  @t  ��  @t  ��   	   1      � $  _�  Y�  _�  @t  !4  @t  !4  Y�   	   1      �   _� �  _�  ��   	   1      � $  _�  ��  _�  �L  �4  �L  �4  ��      1    ,  �� ��  �4 ��  �4 ��  �� ��  �� ��      1    ,  �� q$  �4 q$  �4 ��  �� ��  �� q$      1    ,  !4 q$  .� q$  .� ��  !4 ��  !4 q$      1    ,  !4 ��  0� ��  0� ��  !4 ��  !4 ��      1    ,  y  FP  ��  FP  ��  Y�  y  Y�  y  FP      1    ,  w$  '  ��  '  ��  FP  w$  FP  w$  '      +    ,  �� s  �( s  �( ��  �� ��  �� s      +    ,  �  �  ��  �  ��  #(  �  #(  �  �      +    ,  � ��  �� ��  �� �   � �   � ��      +    ,  @ ��  2� ��  2� ��  @ ��  @ ��      +    ,  @ s  0� s  0� ��  @ ��  @ s      +    ,  �� ��  �( ��  �( ��  �� ��  �� ��      +    ,  w$  HD  ��  HD  ��  W�  w$  W�  w$  HD      +    ,  u0  #(  ��  #(  ��  HD  u0  HD  u0  #(              _�  � GND  +  ,1               _� �8 VDD  +  ,1               <�  � A1 +  ,1               �  � B0 +  ,1               d  � A0 +  ,1               ��  � B1 +  ,1               _�  � Y  +  ,1               _�  � GND               _� �8 VDD               <�  � A1              �  � B0              d  � A0              ��  � B1              _�  � Y      �    , � 	   0  dffs_ni     0    , �4 &� �d &� �d .� �4 .� �4 &�      0    , �4 >\ �d >\ �d F, �4 F, �4 >\      0    , �4 U� �d U� �d ]� �4 ]� �4 U�      1    , � # �| # �| a� � a� � # +  ,1       .    , �� L �� L �� ! �� ! �� L +  ,3       .    , �� w  �� w  �� �� �� �� �� w  +  ,4       .    , �� ! �� ! �� w  �� w  �� !      0    , x� :t q$ :t q$ BD x� BD x� :t      0    , x� Q� q$ Q� q$ Y� x� Y� x� Q�      0    , x� iT q$ iT q$ q$ x� q$ x� iT      1    , |� 6� m< 6� m< u |� u |� 6� +  ,5       .    , iT L a� L a� ! iT ! iT L +  ,6       .    , iT w  a� w  a� �� iT �� iT w  +  ,7       .    , iT ! a� ! a� w  iT w  iT !      0    , Y� &� Q� &� Q� .� Y� .� Y� &�      0    , Y� >\ Q� >\ Q� F, Y� F, Y� >\      0    , Y� U� Q� U� Q� ]� Y� ]� Y� U�      1    , ]� # M� # M� a� ]� a� ]� # +  ,8       +    L L ! L cx Q� cx Q� w  �4 w  �4 cx � cx � ! L !      *    L 4� 	� 4� z� :t z� :t �p �� �p �� z� �� z� �� 	� 4� 	� +  ,10      ,    L D8 @ D8 kH J kH J ~� � ~� � kH �� kH �� @ D8 @      +    < L ! L cx Q� cx Q� w  a� w  a� ! L ! +  ,9       +    < �� ! �� w  �4 w  �4 cx � cx � ! �� ! +  ,2       +    ,  �`  ��  ��  ��  ��  ��  �`  ��  �`  �� +  ,2       0    ,  �<  ��  �  ��  �  ��  �<  ��  �<  ��      0    ,  �<  �4  �  �4  �  �  �<  �  �<  �4      1    ,  �T  ��  ��  ��  ��  ��  �T  ��  �T  �� +  ,1       .    ,  ��  w$ �  w$ �  ��  ��  ��  ��  w$ +  ,3       .    ,  ��  �� �  �� �  ��  ��  ��  ��  �� +  ,4       .    ,  ��  �� �  �� �  ��  ��  ��  ��  ��      0    , |  �� L  �� L  �� |  �� |  ��      0    , |  �4 L  �4 L  � |  � |  �4      1    , �  �� 4  �� 4  �� �  �� �  �� +  ,5       .    ,   w$ &�  w$ &�  ��   ��   w$ +  ,6       .    ,   �� &�  �� &�  ��   ��   �� +  ,7       .    ,   �� &�  �� &�  ��   ��   ��      0    , .�  �� 6�  �� 6�  �� .�  �� .�  ��      0    , .�  �4 6�  �4 6�  � .�  � .�  �4      1    , *�  �� :t  �� :t  �� *�  �� *�  �� +  ,8       +    ,  �`  �� <h  �� <h  ��  �`  ��  �`  ��      )    ,  ��  ix S�  ix S�  �P  ��  �P  ��  ix +  ,10      -    ,  �  y D8  y D8  ��  �  ��  �  y      +    , &�  �� <h  �� <h  �� &�  �� &�  �� +  ,9       0    , 6� &� .� &� .� .� 6� .� 6� &�      0    , 6� >\ .� >\ .� F, 6� F, 6� >\      0    , 6� U� .� U� .� ]� 6� ]� 6� U�      1    , :t # *� # *� a� :t a� :t # +  ,1       .    , &� L  L  ! &� ! &� L +  ,3       .    , &� w   w   �� &� �� &� w  +  ,4       .    , &� !  !  w  &� w  &� !      0    , L :t | :t | BD L BD L :t      0    , L Q� | Q� | Y� L Y� L Q�      0    , L iT | iT | q$ L q$ L iT      1    , 4 6� � 6� � u 4 u 4 6� +  ,5       .    , � L  �� L  �� ! � ! � L +  ,6       .    , � w   �� w   �� �� � �� � w  +  ,7       .    , � !  �� !  �� w  � w  � !      0    ,  � &�  �< &�  �< .�  � .�  � &�      0    ,  � >\  �< >\  �< F,  � F,  � >\      0    ,  � U�  �< U�  �< ]�  � ]�  � U�      1    ,  �� #  �T #  �T a�  �� a�  �� # +  ,8       +    L  �` !  �` cx  �< cx  �< w  6� w  6� cx <h cx <h !  �` !      *    L  �� 	�  �� z�  �� z�  �� �p M� �p M� z� S� z� S� 	�  �� 	� +  ,10      ,    L  � @  � kH  �l kH  �l ~� >\ ~� >\ kH D8 kH D8 @  � @      +    <  �` !  �` cx  �< cx  �< w   �� w   �� !  �` ! +  ,9       +    < &� ! &� w  6� w  6� cx <h cx <h ! &� ! +  ,2       0    ,  L  W�  %  W�  %  _�  L  _�  L  W�      0    ,  L  oT  %  oT  %  w$  L  w$  L  oT      0    ,  L  ��  %  ��  %  ��  L  ��  L  ��      1    ,  d  S�  )  S�  )  �|  d  �|  d  S� +  ,1       .    ,  ,�  HD  4�  HD  4�  R  ,�  R  ,�  HD +  ,3       .    ,  ,�  �p  4�  �p  4�  �4  ,�  �4  ,�  �p +  ,4       .    ,  ,�  R  4�  R  4�  �p  ,�  �p  ,�  R      .    ,  D\  HD  L,  HD  L,  R  D\  R  D\  HD +  ,5       .    ,  D\  �p  L,  �p  L,  �4  D\  �4  D\  �p +  ,6       .    ,  D\  R  L,  R  L,  �p  D\  �p  D\  R      0    ,  S�  W�  [�  W�  [�  _�  S�  _�  S�  W�      0    ,  S�  oT  [�  oT  [�  w$  S�  w$  S�  oT      0    ,  S�  ��  [�  ��  [�  ��  S�  ��  S�  ��      1    ,  P  S�  _�  S�  _�  �|  P  �|  P  S� +  ,7       .    ,  e�  w$  m`  w$  m`  ��  e�  ��  e�  w$ +  ,8       .    ,  e�  �p  m`  �p  m`  �4  e�  �4  e�  �p +  ,9       .    ,  e�  ��  m`  ��  m`  �p  e�  �p  e�  ��      .    ,  }   w$  ��  w$  ��  ��  }   ��  }   w$ +  ,10      .    ,  }   �p  ��  �p  ��  �4  }   �4  }   �p +  ,11      .    ,  }   ��  ��  ��  ��  �p  }   �p  }   ��      0    ,  ��  oT  �d  oT  �d  w$  ��  w$  ��  oT      0    ,  ��  ��  �d  ��  �d  ��  ��  ��  ��  ��      1    ,  ��  kl  �L  kl  �L  �|  ��  �|  ��  kl +  ,12      .    ,  �4  _�  �  _�  �  ix  �4  ix  �4  _� +  ,13      .    ,  �4  �p  �  �p  �  �4  �4  �4  �4  �p +  ,14      .    ,  �4  ix  �  ix  �  �p  �4  �p  �4  ix      .    ,  ��  _�  �t  _�  �t  ix  ��  ix  ��  _� +  ,15      .    ,  ��  �p  �t  �p  �t  �4  ��  �4  ��  �p +  ,16      .    ,  ��  ix  �t  ix  �t  �p  ��  �p  ��  ix      0    ,  �D  oT  �  oT  �  w$  �D  w$  �D  oT      0    ,  �D  ��  �  ��  �  ��  �D  ��  �D  ��      1    ,  �\  kl  ��  kl  ��  �|  �\  �|  �\  kl +  ,17      +    L  a�  R  a�  ��  ��  ��  ��  ix  ��  ix  ��  �p  p  �p  p  R  a�  R      )    <  y  :�  y  R  �`  R  �`  ��      ��      :�  y  :� +  ,19      -    L  ix  J8  ix  y  ��  y  ��  a�  ��  a�  ��  �@  �  �@  �  J8  ix  J8      +    ,  �t  ix  ��  ix  ��  �p  �t  �p  �t  ix +  ,18      +    ,  p  R  ,�  R  ,�  �p  p  �p  p  R +  ,2       +    , �   J8 ؄  J8 ؄  u0 �   u0 �   J8 +  ,2       0    , �$  P �T  P �T  W� �$  W� �$  P      0    , �$  g� �T  g� �T  oT �$  oT �$  g�      1    , �  L, �l  L, �l  s< �  s< �  L, +  ,1       .    , ؄  @t д  @t д  J8 ؄  J8 ؄  @t +  ,3       .    , ؄  u0 д  u0 д  ~� ؄  ~� ؄  u0 +  ,4       .    , ؄  J8 д  J8 д  u0 ؄  u0 ؄  J8      0    , ��  P �  P �  W� ��  W� ��  P      0    , ��  g� �  g� �  oT ��  oT ��  g�      1    , ��  L, �,  L, �,  s< ��  s< ��  L, +  ,5       .    , �D  @t �t  @t �t  J8 �D  J8 �D  @t +  ,6       .    , �D  u0 �t  u0 �t  ~� �D  ~� �D  u0 +  ,7       .    , �D  J8 �t  J8 �t  u0 �D  u0 �D  J8      0    , ��  P ��  P ��  W� ��  W� ��  P      0    , ��  g� ��  g� ��  oT ��  oT ��  g�      1    , ��  L, ��  L, ��  s< ��  s< ��  L, +  ,8       +    , �   J8 ��  J8 ��  u0 �   u0 �   J8      )    , p  2� ��  2� ��  �� p  �� p  2� +  ,10      -    , ��  Bh �(  Bh �(  }  ��  }  ��  Bh      +    , �t  J8 ��  J8 ��  u0 �t  u0 �t  J8 +  ,9       +    , L  �� a�  �� a�  �� L  �� L  �� +  ,2       0    , Q�  �� Y�  �� Y�  �� Q�  �� Q�  ��      0    , Q�  �4 Y�  �4 Y�  � Q�  � Q�  �4      1    , M�  �� ]�  �� ]�  �� M�  �� M�  �� +  ,1       .    , a�  w$ iT  w$ iT  �� a�  �� a�  w$ +  ,3       .    , a�  �� iT  �� iT  �� a�  �� a�  �� +  ,4       .    , a�  �� iT  �� iT  �� a�  �� a�  ��      0    , q$  �� x�  �� x�  �� q$  �� q$  ��      0    , q$  �4 x�  �4 x�  � q$  � q$  �4      1    , m<  �� |�  �� |�  �� m<  �� m<  �� +  ,5       .    , ��  w$ ��  w$ ��  �� ��  �� ��  w$ +  ,6       .    , ��  �� ��  �� ��  �� ��  �� ��  �� +  ,7       .    , ��  �� ��  �� ��  �� ��  �� ��  ��      0    , �d  �� �4  �� �4  �� �d  �� �d  ��      0    , �d  �4 �4  �4 �4  � �d  � �d  �4      1    , �|  �� �  �� �  �� �|  �� �|  �� +  ,8       +    , L  �� �  �� �  �� L  �� L  ��      )    , 4�  ix ��  ix ��  �P 4�  �P 4�  ix +  ,10      -    , D8  y ��  y ��  �� D8  �� D8  y      +    , ��  �� �  �� �  �� ��  �� ��  �� +  ,9       0    , �   �| ��  �| ��  �L �   �L �   �|      1    , �8  �� ��  �� ��  �4 �8  �4 �8  �� +  ,1       .    , ��  �� ܐ  �� ܐ  �� ��  �� ��  �� +  ,3       .    , ��  �( ܐ  �( ܐ  �� ��  �� ��  �( +  ,4       .    , ��  �� ܐ  �� ܐ  �( ��  �( ��  ��      0    , �T  c� �$  c� �$  kl �T  kl �T  c�      0    , �T  { �$  { �$  �� �T  �� �T  {      0    , �T  �| �$  �| �$  �L �T  �L �T  �|      1    , �l  _� �  _� �  �4 �l  �4 �l  _� +  ,5       .    , ��  S� ��  S� ��  ]� ��  ]� ��  S� +  ,6       .    , ��  �( ��  �( ��  �� ��  �� ��  �( +  ,7       .    , ��  ]� ��  ]� ��  �( ��  �( ��  ]�      .    , d  S� 4  S� 4  ]� d  ]� d  S� +  ,8       .    , d  �( 4  �( 4  �� d  �� d  �( +  ,9       .    , d  ]� 4  ]� 4  �( d  �( d  ]�      0    ,   c� $�  c� $�  kl   kl   c�      0    ,   { $�  { $�  ��   ��   {      0    ,   �| $�  �| $�  �L   �L   �|      1    ,   _� (�  _� (�  �4   �4   _� +  ,10      .    , .�  �� 6h  �� 6h  �� .�  �� .�  �� +  ,11      .    , .�  �( 6h  �( 6h  �� .�  �� .�  �( +  ,12      .    , .�  �� 6h  �� 6h  �( .�  �( .�  ��      .    , F  �� M�  �� M�  �� F  �� F  �� +  ,13      .    , F  �( M�  �( M�  �� F  �� F  �( +  ,14      .    , F  �� M�  �� M�  �( F  �( F  ��      0    , U�  �| ]x  �| ]x  �L U�  �L U�  �|      1    , Q�  �� a`  �� a`  �4 Q�  �4 Q�  �� +  ,15      +    L *�  ]� *�  �� cT  �� cT  �( �D  �( �D  �� �x  �� �x  ]� *�  ]�      )    L B   FP B   u0 z�  u0 z�  �� ��  �� ��  u0 �  u0 �  FP B   FP +  ,17      -    L 2�  U� 2�  �� k$  �� k$  �� �t  �� �t  �� ب  �� ب  U� 2�  U�      +    , M�  �� cT  �� cT  �( M�  �( M�  �� +  ,16      +    , �D  �� ��  �� ��  �( �D  �( �D  �� +  ,2       +    , Y�  J8 o  J8 o  ]� Y�  ]� Y�  J8 +  ,2       0    , _l  P g<  P g<  W� _l  W� _l  P      1    , [�  L, k$  L, k$  [� [�  [� [�  L, +  ,1       .    , o  @t v�  @t v�  J8 o  J8 o  @t +  ,3       .    , o  ]� v�  ]� v�  g� o  g� o  ]� +  ,4       .    , o  J8 v�  J8 v�  ]� o  ]� o  J8      0    , ~�  P �|  P �|  W� ~�  W� ~�  P      1    , z�  L, �d  L, �d  [� z�  [� z�  L, +  ,5       +    , Y�  J8 �X  J8 �X  ]� Y�  ]� Y�  J8      )    , B   2� ��  2� ��  u0 B   u0 B   2� +  ,7       -    , Q�  Bh �(  Bh �(  e� Q�  e� Q�  Bh      +    , v�  J8 �X  J8 �X  ]� v�  ]� v�  J8 +  ,6       0    ,  L   %   % &�  L &�  L       0    ,  L 6�  % 6�  % >\  L >\  L 6�      0    ,  L M�  % M�  % U�  L U�  L M�      0    ,  L el  % el  % m<  L m<  L el      0    ,  L |�  % |�  % ��  L ��  L |�      1    ,  d 4  ) 4  ) ��  d ��  d 4 +  ,1       .    ,  ,� �  4� �  4� �  ,� �  ,� � +  ,3       .    ,  ,� ��  4� ��  4� �L  ,� �L  ,� �� +  ,4       .    ,  ,� �  4� �  4� ��  ,� ��  ,� �      .    ,  D\ �  L, �  L, �  D\ �  D\ � +  ,5       .    ,  D\ ��  L, ��  L, �L  D\ �L  D\ �� +  ,6       .    ,  D\ �  L, �  L, ��  D\ ��  D\ �      0    ,  S� d  [� d  [� 4  S� 4  S� d      0    ,  S� *�  [� *�  [� 2�  S� 2�  S� *�      0    ,  S� BD  [� BD  [� J  S� J  S� BD      0    ,  S� Y�  [� Y�  [� a�  S� a�  S� Y�      0    ,  S� q$  [� q$  [� x�  S� x�  S� q$      1    ,  P |  _� |  _� |�  P |�  P | +  ,7       .    ,  e� W�  m` W�  m` a�  e� a�  e� W� +  ,8       .    ,  e� u  m` u  m` ~�  e� ~�  e� u +  ,9       .    ,  e� a�  m` a�  m` u  e� u  e� a�      .    ,  }  W�  �� W�  �� a�  }  a�  }  W� +  ,10      .    ,  }  u  �� u  �� ~�  }  ~�  }  u +  ,11      .    ,  }  a�  �� a�  �� u  }  u  }  a�      0    ,  �� O�  �d O�  �d W�  �� W�  �� O�      0    ,  �� g`  �d g`  �d o0  �� o0  �� g`      1    ,  �� L  �L L  �L s  �� s  �� L +  ,12      .    ,  �4 0�  � 0�  � :t  �4 :t  �4 0� +  ,13      .    ,  �4 u  � u  � ~�  �4 ~�  �4 u +  ,14      .    ,  �4 :t  � :t  � u  �4 u  �4 :t      0    ,  �� @P  �� @P  �� H   �� H   �� @P      0    ,  �� W�  �� W�  �� _�  �� _�  �� W�      1    ,  �� <h  �� <h  �� cx  �� cx  �� <h +  ,15      .    ,  �t 0�  �D 0�  �D :t  �t :t  �t 0� +  ,16      .    ,  �t u  �D u  �D ~�  �t ~�  �t u +  ,17      .    ,  �t :t  �D :t  �D u  �t u  �t :t      0    ,  � O�  �� O�  �� W�  � W�  � O�      0    ,  � g`  �� g`  �� o0  � o0  � g`      1    ,  �, L  �� L  �� s  �, s  �, L +  ,18      +    �  a� �  a� a�  �� a�  �� J  �� J  �� :t  �� :t  �� J  �� J  �� u  a� u  a� ~�  [� ~�  [� ��  p ��  p @  L @  L �  a� �      *    |  y  �  y #  �T #  �T 2�  �0 2�  �0 �|  y �|  y �@  s< �@  s< ��     ��     �  � �  �  �  y  � +  ,20      ,    �  ix �  ix Y�  �� Y�  �� BD  �� BD  �� 2�  ܴ 2�  ܴ BD  � BD  � |�  ix |�  ix ��  c� ��  c� �X  � �X  � p  | p  | �  ix �      +    <  �� :t  �� J  �� J  �� u  �D u  �D :t  �� :t +  ,19      +    <  ,� �  ,� ��  p ��  p @  L @  L �  ,� � +  ,2       0    , �$ :t �T :t �T BD �$ BD �$ :t      0    , �$ Q� �T Q� �T Y� �$ Y� �$ Q�      0    , �$ iT �T iT �T q$ �$ q$ �$ iT      1    , � 6� �l 6� �l u � u � 6� +  ,1       .    , ؄ *� д *� д 4� ؄ 4� ؄ *� +  ,3       .    , ؄ �� д �� д �L ؄ �L ؄ �� +  ,4       .    , ؄ 4� д 4� д �� ؄ �� ؄ 4�      0    , �� M� � M� � U� �� U� �� M�      0    , �� el � el � m< �� m< �� el      0    , �� |� � |� � �� �� �� �� |�      1    , �� J �, J �, �� �� �� �� J +  ,5       .    , �D *� �t *� �t 4� �D 4� �D *� +  ,6       .    , �D �� �t �� �t �L �D �L �D �� +  ,7       .    , �D 4� �t 4� �t �� �D �� �D 4�      0    , �� :t �� :t �� BD �� BD �� :t      0    , �� Q� �� Q� �� Y� �� Y� �� Q�      0    , �� iT �� iT �� q$ �� q$ �� iT      1    , �� 6� �� 6� �� u �� u �� 6� +  ,8       +    L �� 4� �� w  �� w  �� �� �$ �� �$ w  �  w  �  4� �� 4�      *    L �� ( �� �p �d �p �d �� �� �� �� �p p �p p ( �� ( +  ,10      ,    L �( ,� �( ~� � ~� � �X �� �X �� ~� �� ~� �� ,� �( ,�      +    < �� 4� �� w  �� w  �� �� �t �� �t 4� �� 4� +  ,9       +    < ؄ 4� ؄ �� �$ �� �$ w  �  w  �  4� ؄ 4� +  ,2       0    , �  d �� d �� 4 �  4 �  d      1    , �8 | �� | ��  �8  �8 | +  ,1       .    , �� � ܐ � ܐ � �� � �� � +  ,3       .    , �� ! ܐ ! ܐ *� �� *� �� ! +  ,4       .    , �� � ܐ � ܐ ! �� ! �� �      0    , �T  �$  �$ &� �T &� �T       0    , �T 6� �$ 6� �$ >\ �T >\ �T 6�      0    , �T M� �$ M� �$ U� �T U� �T M�      0    , �T el �$ el �$ m< �T m< �T el      0    , �T |� �$ |� �$ �� �T �� �T |�      1    , �l 4 � 4 � �� �l �� �l 4 +  ,5       .    , �� � �� � �� � �� � �� � +  ,6       .    , �� �� �� �� �� �L �� �L �� �� +  ,7       .    , �� � �� � �� �� �� �� �� �      .    , d � 4 � 4 � d � d � +  ,8       .    , d �� 4 �� 4 �L d �L d �� +  ,9       .    , d � 4 � 4 �� d �� d �      0    ,   $�  $� &�  &�        0    ,  6� $� 6� $� >\  >\  6�      0    ,  M� $� M� $� U�  U�  M�      0    ,  el $� el $� m<  m<  el      0    ,  |� $� |� $� ��  ��  |�      1    ,  4 (� 4 (� ��  ��  4 +  ,10      .    , .� *� 6h *� 6h 4� .� 4� .� *� +  ,11      .    , .� H  6h H  6h Q� .� Q� .� H  +  ,12      .    , .� 4� 6h 4� 6h H  .� H  .� 4�      0    , >8 :t F :t F BD >8 BD >8 :t      1    , :P 6� I� 6� I� F, :P F, :P 6� +  ,13      .    , M� *� U� *� U� 4� M� 4� M� *� +  ,14      .    , M� H  U� H  U� Q� M� Q� M� H  +  ,15      .    , M� 4� U� 4� U� H  M� H  M� 4�      0    , _l # g< # g< *� _l *� _l #      0    , _l :t g< :t g< BD _l BD _l :t      1    , [�  k$  k$ F, [� F, [�  +  ,16      .    , o d v� d v� ( o ( o d +  ,17      .    , o H  v� H  v� Q� o Q� o H  +  ,18      .    , o ( v� ( v� H  o H  o (      0    , ~� # �| # �| *� ~� *� ~� #      0    , ~� :t �| :t �| BD ~� BD ~� :t      1    , z�  �d  �d F, z� F, z�  +  ,19      +    | $� � $� @ *� @ *� 4� Y� 4� Y� ( �X ( �X H  *� H  *� �� �x �� �x ! �D ! �D � $� �      *    l <D  � <D � B  � B  � �� � �� _� B  _� B  �� � �� � 8� �� 8� ��  � <D  � +  ,21      ,    | ,� � ,� p 2� p 2� ,� Q� ,� Q� X �( X �( O� 2� O� 2� �X ب �X ب (� �t (� �t � ,� �      +    , v� ( �X ( �X H  v� H  v� ( +  ,20      +    , �D � �� � �� ! �D ! �D � +  ,2    
  via  �  B�        m<  �   
  via  �  B�        ��  �   
  via  �  B�         Bh  �   
  via  �  B�        �  �   
  via  �  B�        �$  �      1    ,         p     p  '      '              1    ,     �� p �� p ��     ��     ��      3    , �  �P X  �P X  �� �  �� �  �P      3    , cx  �P w   �P w   �� cx  �� cx  �P      3    ,  8�  �P  L,  �P  L,  ��  8�  ��  8�  �P      3    , �`  �P ��  �P ��  �� �`  �� �`  �P      3    , �  �P ��  �P ��  �� �  �� �  �P      -    ,  ~�  a�  ��  a�  ��  y  ~�  y  ~�  a�      /    , 8�  ix @P  ix @P  qH 8�  qH 8�  ix      /    ,  �$  HD  ��  HD  ��  P  �$  P  �$  HD      /    ,  �D  D\  �  D\  �  L,  �D  L,  �D  D\      /    , Q�  6� Y�  6� Y�  >� Q�  >� Q�  6�      /    , �d  D\ �4  D\ �4  L, �d  L, �d  D\      1    , 4�  e� D8  e� D8  u0 4�  u0 4�  e�      1    ,  p  '  '  '  '  @t  p  @t  p  '      1    ,  d  @t  '  @t  '  S�  d  S�  d  @t   	   1      �   �|  P  �|  '      1    ,  ��  _�  �X  _�  �X  kl  ��  kl  ��  _�      1    ,  ��  P  �X  P  �X  _�  ��  _�  ��  P      1    , �   8� ��  8� ��  L, �   L, �   8�      1    , �,  ' ��  ' ��  8� �,  8� �,  '      1    , [�  8� i0  8� i0  L, [�  L, [�  8�      1    , Y�  ' i0  ' i0  8� Y�  8� Y�  '   	   1      �  "�  >� "�  '      1    ,   N  (�  N  (�  _�   _�   N       1    ,   >� *�  >� *�  N    N    >�      1    ,  �<  D\  ��  D\  ��  S�  �<  S�  �<  D\   	   1      �   �,  kl  �,  P      1    , M�  2� ]�  2� ]�  Bh M�  Bh M�  2�      1    ,  �\  @t  ��  @t  ��  P  �\  P  �\  @t      1    , �|  @t �  @t �  P �|  P �|  @t      +    ,   <� ,�  <� ,�  P   P   <�      +    ,  |  #(  )  #(  )  Bh  |  Bh  |  #(      +    ,  p  Bh  )  Bh  )  R  p  R  p  Bh      +    ,  ��  a�  �L  a�  �L  ix  ��  ix  ��  a�      +    ,  ��  N   �L  N   �L  a�  ��  a�  ��  N       +    , �,  :� ��  :� ��  J8 �,  J8 �,  :�      +    , �8  #( ��  #( ��  :� �8  :� �8  #(      +    , Y�  :� k$  :� k$  J8 Y�  J8 Y�  :�      +    , W�  #( k$  #( k$  :� W�  :� W�  #(      +    ,   P *�  P *�  ]�   ]�   P      +    ,  |  � �  � �  #(  |  #(  |  �      ,    , L  *� 4t  *� 4t  U� L  U� L  *�      ,    ,  �  *�  0�  *�  0�  J8  �  J8  �  *�      ,    ,  ~�  FP  �  FP  �  a�  ~�  a�  ~�  FP      ,    , �h  *� ֐  *� ֐  Bh �h  Bh �h  *�      ,    , O�  *� r�  *� r�  Bh O�  Bh O�  *�      ,    ,  �  � ��  � ��  *�  �  *�  �  �      0    , �  Bh &�  Bh &�  J8 �  J8 �  Bh      0    , �L  | �  | �  L �L  L �L  |      0    , |�  | ��  | ��  L |�  L |�  |      0    , el  | m<  | m<  L el  L el  |      0    , M�  | U�  | U�  L M�  L M�  |      0    , 6�  | >\  | >\  L 6�  L 6�  |      0    ,   | &�  | &�  L   L   |      0    , �  | |  | |  L �  L �  |      0    ,  �<  |  �  |  �  L  �<  L  �<  |      0    ,  ��  |  ��  |  ��  L  ��  L  ��  |      0    ,  �\  |  �,  |  �,  L  �\  L  �\  |      0    ,  ��  |  ��  |  ��  L  ��  L  ��  |      0    ,  �|  |  �L  |  �L  L  �|  L  �|  |      0    ,  {  |  ��  |  ��  L  {  L  {  |      0    ,  c�  |  kl  |  kl  L  c�  L  c�  |      0    ,  L,  |  S�  |  S�  L  L,  L  L,  |      0    ,  4�  |  <�  |  <�  L  4�  L  4�  |      0    ,  L  |  %  |  %  L  L  L  L  |      0    ,  X  0�  #(  0�  #(  8�  X  8�  X  0�      0    ,  ��  S�  �p  S�  �p  [�  ��  [�  ��  S�      0    , �  ,� ��  ,� ��  4� �  4� �  ,�      0    , ]x  ,� eH  ,� eH  4� ]x  4� ]x  ,�      0    , ��  | ��  | ��  L ��  L ��  |      0    , �,  | ��  | ��  L �,  L �,  |      0    , ڜ  | �l  | �l  L ڜ  L ڜ  |      0    , �  | ��  | ��  L �  L �  |      0    , 	|  | L  | L  L 	|  L 	|  |      0    ,  �  | (�  | (�  L  �  L  �  |      0    , 8\  | @,  | @,  L 8\  L 8\  |      0    , O�  | W�  | W�  L O�  L O�  |      0    , g<  | o  | o  L g<  L g<  |      0    , ~�  | �|  | �|  L ~�  L ~�  |      0    , �  | ��  | ��  L �  L �  |      0    , ��  | �\  | �\  L ��  L ��  |      0    , ��  | ��  | ��  L ��  L ��  |      0    , �l  | �<  | �<  L �l  L �l  |             ��  � GND  +  ,1       .    , 2�  c� F,  c� F,  w$ 2�  w$ 2�  c�      .    ,  �H  Bh �  Bh �  U�  �H  U�  �H  Bh   	   .      � , #  w$ #  g�  ��  g�  ��  N   ��  N    	   .      �   ix  w$  ix  Bh  �h  Bh      .    ,  �h  >�  ��  >�  ��  R  �h  R  �h  >�      .    , L  0� _�  0� _�  D\ L  D\ L  0�   	   .      �   0�  HD  0�  .� _�  .�   	   .      �  L  S� L  Bh �  Bh      .    , ��  >� �  >� �  R ��  R ��  >�   	   .      � $ F,  g� ��  g� ��  U� ��  U�      0    ,  L �t  % �t  % �D  L �D  L �t      0    , �l �t �< �t �< �D �l �D �l �t      0    , �� �t �� �t �� �D �� �D �� �t      0    , �� �t �\ �t �\ �D �� �D �� �t      0    , � �t �� �t �� �D � �D � �t      0    , ~� �t �| �t �| �D ~� �D ~� �t      0    , g< �t o �t o �D g< �D g< �t      0    , O� �t W� �t W� �D O� �D O� �t      0    , 8\ �t @, �t @, �D 8\ �D 8\ �t      0    ,  � �t (� �t (� �D  � �D  � �t      0    , 	| �t L �t L �D 	| �D 	| �t      0    , � �t �� �t �� �D � �D � �t      0    , ڜ �t �l �t �l �D ڜ �D ڜ �t      0    , �, �t �� �t �� �D �, �D �, �t      0    , �� �t �� �t �� �D �� �D �� �t      0    , �L �t � �t � �D �L �D �L �t      0    , |� �t �� �t �� �D |� �D |� �t      0    , el �t m< �t m< �D el �D el �t      0    , M� �t U� �t U� �D M� �D M� �t      0    , 6� �t >\ �t >\ �D 6� �D 6� �t      0    ,  �t &� �t &� �D  �D  �t      0    , � �t | �t | �D � �D � �t      0    ,  �< �t  � �t  � �D  �< �D  �< �t      0    ,  �� �t  �� �t  �� �D  �� �D  �� �t      0    ,  �\ �t  �, �t  �, �D  �\ �D  �\ �t      0    ,  �� �t  �� �t  �� �D  �� �D  �� �t      0    ,  �| �t  �L �t  �L �D  �| �D  �| �t      0    ,  { �t  �� �t  �� �D  { �D  { �t      0    ,  c� �t  kl �t  kl �D  c� �D  c� �t      0    ,  L, �t  S� �t  S� �D  L, �D  L, �t      0    ,  4� �t  <� �t  <� �D  4� �D  4� �t      0    , ]x ]� eH ]� eH el ]x el ]x ]�      0    , 8\ el @, el @, m< 8\ m< 8\ el      0    , 8\ |� @, |� @, �� 8\ �� 8\ |�      0    , � � �� � �� �� � �� � �      0    ,  X �  #( �  #( ��  X ��  X �      0    , q$ �| x� �| x� �L q$ �L q$ �|      +    ,  | �� � �� � �   | �   | ��      +    , Y� H  k$ H  k$ W� Y� W� Y� H       +    , W� W� k$ W� k$ kH W� kH W� W�      +    , �8 �( �� �( �� �� �8 �� �8 �(      +    , *� _� F _� F �� *� �� *� _�      +    , �, �� �� �� �� �( �, �( �, ��      +    ,  | �(  ) �(  ) ��  | ��  | �(      +    ,  p ��  ) ��  ) �(  p �(  p ��      +    , m< w  |� w  |� �� m< �� m< w       +    , kH �� ~� �� ~� �( kH �( kH ��      /    , g`  �, o0  �, o0  �� g`  �� g`  �,      /    ,  >�  �,  FP  �,  FP  ��  >�  ��  >�  �,      /    , �  �, �  �, �  �� �  �� �  �,      /    ,  �D �  � �  � d  �D d  �D �      /    , ڜ �@ �l �@ �l � ڜ � ڜ �@      /    , �� � Ҩ � Ҩ | �� | �� �      /    , 2�  ܴ :P  ܴ :P  � 2�  � 2�  ܴ      /    , L  ܴ   ܴ   � L  � L  ܴ      /    , ܐ  ܴ �`  ܴ �`  � ܐ  � ܐ  ܴ      /    , z�  �0 ��  �0 ��  �  z�  �  z�  �0      /    , �� M� �t M� �t U� �� U� �� M�      /    , H  �� O� �� O� �d H  �d H  ��      /    , �p �@ �@ �@ �@ � �p � �p �@      /    ,  '  �  .�  �  .�  ��  '  ��  '  �      /    ,  qH 4�  y 4�  y <h  qH <h  qH 4�      /    ,  ��  �,  �X  �,  �X  ��  ��  ��  ��  �,      /    ,  _�  �x  g�  �x  g�  �H  _�  �H  _�  �x      1    , Y� Y� i0 Y� i0 iT Y� iT Y� Y�      1    , cx  �D s  �D s  �� cx  �� cx  �D      1    ,  :�  �D  J8  �D  J8  ��  :�  ��  :�  �D      1    , �  �D p  �D p  �� �  �� �  �D   	   1      �   �` |  �� |      1    ,  �\ �  �� �  �� L  �\ L  �\ �   	   1      �   �<  �4  �< .�   	   1      �  6�  �4 6� .�      1    , �� � ֐ � ֐ d �� d �� �   	   1      �  �� BD ��  g�   	   1      �  �$  g� �$ BD   	   1      �  �� � �� �      1    , ִ �X �T �X �T �� ִ �� ִ �X   	   1      �  �x �X �x �� �l ��      1    , [� F, i0 F, i0 Y� [� Y� [� F,      1    , �, � �� � �� �� �, �� �, �      1    , �  �� �� �� �� � �  � �  ��   	   1      �  cT iT cT ��      1    , (� a� D a� D �� (� �� (� a�   	   1      �   � ��  � ��      1    ,  p �  ' �  ' ��  p ��  p �      1    ,  d ��  ' ��  ' �  d �  d ��   	   1      �   �� s  �� ��   	   1      �   �| s  �| ��   	   1      �  ��  ��  [�   	   1      �  |�  �� >8  ��   	   1      � $ �� | �� � @, � @, 6�      1    , .�  �� >8  �� >8  �l .�  �l .�  ��   	   1      � $ ��  �4 ��  �� W�  �� W�  �4   	   1      � $ �l 4� �� 4� ��  y �l  y   	   1      �  � | �  �4   	   1      �  d  �� �H  ��   	   1      �  Q�  �4 Q� .�   	   1      �  w   � W�  �   	   1      �  �4  �4 �4 .�      1    , d  ��   ��   �l d  �l d  ��      1    , ب  �� �H  �� �H  �l ب  �l ب  ��      1    , w   �H ��  �H ��  �� w   �� w   �H   	   1      �  d u d ��   	   1      �  �� Q� � Q�   	   1      �  S� a� S� �L   	   1      �  u �4 u ��   	   1      �  �L a� �L �(      1    , �� J �\ J �\ Y� �� Y� �� J      1    , D8 �� S� �� S� �L D8 �L D8 ��      1    , �� �X �( �X �( �� �� �� �� �X      1    , o0 u z� u z� �� o0 �� o0 u      1    , m< �� |� �� |� �4 m< �4 m< ��   	   1      �   }  6�  �� 6�   	   1      � $  �� 0�  ��  �  �8  �  �8  �|   	   1      � ,  _� X  �� X  ��  ��  W�  ��  W�  �|   	   1      �   [�  �T  ,�  �T  ,�  �$      1    ,  #(  �$  2�  �$  2� �  #( �  #(  �$      1    ,  m` 0�  }  0�  }  @P  m` @P  m` 0�      1    ,  ��  �D  �@  �D  �@  ��  ��  ��  ��  �D      1    ,  [�  �  kl  �  kl  �0  [�  �0  [�  �   	   1      �  u  �� u  '   	   1      �   �  ��  �  S�   	   1      �  d  �� d  '   	   1      �  U�  �� U�  Bh   	   1      �  �L  P �L  ��   	   1      �  4�  �� 4�  e�      *    ,      � p  � p ��     ��      �      )    ,         p     p  �P      �P                     �  � S  +  ,1              m<  � CLK  +  ,1               Bh  � D  +  ,1              �$  � Q  +  ,1              ��  � QB +  ,1              �� �8 VDD  +  ,1       .    , a�  �P u  �P u  �� a�  �� a�  �P      .    ,  8�  �P  L,  �P  L,  ��  8�  ��  8�  �P      .    ,  ��  �P d  �P d  ��  ��  ��  ��  �P      .    ,  �h �  �� �  �� @  �h @  �h �   	   .      � $  �\ 0�  �\  ��  ��  ��  ��  �4   	   .      � $ �t &� �( &� �( U� v� U�   	   .      �  Ԝ *� Ԝ  ~�   	   .      � < �  R (�  R (�  S� u  S� u  .� I�  .� I�  ��   	   .      �  �\  ~� �\ *�      .    , �� �d �H �d �H �� �� �� �� �d      .    , �� � ؄ � ؄ X �� X �� �   	   .      �  r�  g� r� d   	   .      � $ Q� *� Q�  �t I�  �t I�  ��   	   .      �  2� *� 2�  ��      .    , ,�  �� @,  �� @,  �` ,�  �` ,�  ��   	   .      �  ��  �� �� �   	   .      �  L � L  �`   	   .      �  ب  �� ب  �`   	   .      �  ��  �x ��  �x   	   .      �  el L el  ��   	   .      �  ��  �� �� L      .    , p  �� �  �� �  �` p  �` p  ��      .    , ִ  �� �<  �� �<  �` ִ  �` ִ  ��      .    , u  �T ��  �T ��  �� u  �� u  �T   	   .      �  ب *� ب L �P L      .    , �� H  �P H  �P [� �� [� �� H       .    , BD �� U� �� U� �@ BD �@ BD ��      .    , �� �d � �d � �� �� �� �� �d   	   .      �   ix W�  ix .�   	   .      �   �  �4  � 0�   	   .      � $  ��  �4  ��  ��  ix  ��  ix  ��   	   .      �   HD �  HD  �4      .    ,  !4  �0  4�  �0  4� �  !4 �  !4  �0      .    ,  kl .�  ~� .�  ~� BD  kl BD  kl .�      .    ,  ��  �P  �4  �P  �4  ��  ��  ��  ��  �P      .    ,  Y�  ��  m`  ��  m`  �$  Y�  �$  Y�  ��   	   .      �  BD �X  �� �X  �� ~�   	   .      �   0� �L  0� �� � ��   	   .      �  � L �  ��   	   .      �  #  �� # L   	   .      �  �� �� r� �� r� Q�      -    ,  � �� �� �� �� ��  � ��  � ��      -    , M� O� r� O� r� s M� s M� O�      -    , 2� O� M� O� M� �X 2� �X 2� O�      -    , �h �X ֐ �X ֐ �� �h �� �h �X      -    ,  � �X  0� �X  0� ��  � ��  � �X      -    , cx ~� �� ~� �� �� cx �� cx ~�      -    ,  ��  y  �  y  �  �@  ��  �@  ��  y             �  � S              m<  � CLK               Bh  � D              �$  � Q              ��  � QB             ��  � GND              �� �8 VDD      �     � 	   1  or03    +    ,  p  J8  ,�  J8  ,�  ]�  p  ]�  p  J8 +  ,2       0    ,  L  P  %  P  %  W�  L  W�  L  P      1    ,  d  L,  )  L,  )  [�  d  [�  d  L, +  ,1       .    ,  ,�  @t  4�  @t  4�  J8  ,�  J8  ,�  @t +  ,3       .    ,  ,�  ]�  4�  ]�  4�  g�  ,�  g�  ,�  ]� +  ,4       .    ,  ,�  J8  4�  J8  4�  ]�  ,�  ]�  ,�  J8      0    ,  <�  P  D\  P  D\  W�  <�  W�  <�  P      1    ,  8�  L,  HD  L,  HD  [�  8�  [�  8�  L, +  ,5       .    ,  L,  @t  S�  @t  S�  J8  L,  J8  L,  @t +  ,6       .    ,  L,  a�  S�  a�  S�  kl  L,  kl  L,  a� +  ,7       .    ,  L,  J8  S�  J8  S�  a�  L,  a�  L,  J8      0    ,  [�  S�  c�  S�  c�  [�  [�  [�  [�  S�      1    ,  W�  P  g�  P  g�  _�  W�  _�  W�  P +  ,8       .    ,  kl  @t  s<  @t  s<  J8  kl  J8  kl  @t +  ,9       .    ,  kl  a�  s<  a�  s<  kl  kl  kl  kl  a� +  ,10      .    ,  kl  J8  s<  J8  s<  a�  kl  a�  kl  J8      0    ,  {  P  ��  P  ��  W�  {  W�  {  P      1    ,  w$  L,  ��  L,  ��  [�  w$  [�  w$  L, +  ,11      .    ,  ��  @t  �|  @t  �|  J8  ��  J8  ��  @t +  ,12      .    ,  ��  a�  �|  a�  �|  kl  ��  kl  ��  a� +  ,13      .    ,  ��  J8  �|  J8  �|  a�  ��  a�  ��  J8      0    ,  �L  S�  �  S�  �  [�  �L  [�  �L  S�      1    ,  �d  P  �  P  �  _�  �d  _�  �d  P +  ,14      +    L  �  J8  �  N   ��  N   ��  a�  <�  a�  <�  ]�  p  ]�  p  J8  �  J8      )    L  ��  2�  ��  6�  �h  6�  �h  y  %  y  %  u0      u0      2�  ��  2� +  ,16      -    L  ��  Bh  ��  FP  ��  FP  ��  ix  4�  ix  4�  e�  �  e�  �  Bh  ��  Bh      +    <  �  J8  �  N   ��  N   ��  a�  �|  a�  �|  J8  �  J8 +  ,15      0    ,  L d  % d  % 4  L 4  L d      0    ,  L *�  % *�  % 2�  L 2�  L *�      1    ,  d |  ) |  ) 6�  d 6�  d | +  ,1       .    ,  ,� �  4� �  4� �  ,� �  ,� � +  ,3       .    ,  ,� 8�  4� 8�  4� BD  ,� BD  ,� 8� +  ,4       .    ,  ,� �  4� �  4� 8�  ,� 8�  ,� �      0    ,  >�   FP   FP &�  >� &�  >�       0    ,  >� 6�  FP 6�  FP >\  >� >\  >� 6�      0    ,  >� M�  FP M�  FP U�  >� U�  >� M�      0    ,  >� el  FP el  FP m<  >� m<  >� el      0    ,  >� |�  FP |�  FP ��  >� ��  >� |�      1    ,  :� 4  J8 4  J8 ��  :� ��  :� 4 +  ,5       .    ,  N  �  U� �  U� �  N  �  N  � +  ,6       .    ,  N  ��  U� ��  U� �L  N  �L  N  �� +  ,7       .    ,  N  �  U� �  U� ��  N  ��  N  �      .    ,  e� �  m` �  m` �  e� �  e� � +  ,8       .    ,  e� ��  m` ��  m` �L  e� �L  e� �� +  ,9       .    ,  e� �  m` �  m` ��  e� ��  e� �      .    ,  }  �  �� �  �� �  }  �  }  � +  ,10      .    ,  }  ��  �� ��  �� �L  }  �L  }  �� +  ,11      .    ,  }  �  �� �  �� ��  }  ��  }  �      0    ,  �� d  �p d  �p 4  �� 4  �� d      0    ,  �� *�  �p *�  �p 2�  �� 2�  �� *�      0    ,  �� BD  �p BD  �p J  �� J  �� BD      0    ,  �� Y�  �p Y�  �p a�  �� a�  �� Y�      0    ,  �� q$  �p q$  �p x�  �� x�  �� q$      1    ,  �� |  �X |  �X |�  �� |�  �� | +  ,12      +    L  �L �  �L ~�  �p ~�  �p ��  8� ��  8� 8�  p 8�  p �  �L �      *    L  ��  �  �� �@  �� �@  �� ��  !4 ��  !4 O�     O�      �  ��  � +  ,14      ,    L  � �  � ��  �@ ��  �@ �X  0� �X  0� @P  � @P  � �  � �      +    <  �L �  �L ~�  �p ~�  �p ��  �� ��  �� �  �L � +  ,13      +    ,  p �  ,� �  ,� 8�  p 8�  p � +  ,2    
  via    oT  ��   
  via    �|  ��   
  via    L,  ��   
  via    L  ��      1    ,     ��  �h ��  �h ��     ��     ��      1    ,          �h      �h  '      '              3    ,  ��  ��  �@  ��  �@  �P  ��  �P  ��  ��      3    ,  e�  ��  y  ��  y  �P  e�  �P  e�  ��      3    ,  Bh  ��  U�  ��  U�  �P  Bh  �P  Bh  ��      3    ,  �  ��  '  ��  '  �P  �  �P  �  ��      �    ,          �h      �h ��     ��              )    ,          �h      �h  y      y              *    ,      �  �h  �  �h ��     ��      �      ,    ,  m`  *�  ��  *�  ��  Bh  m`  Bh  m`  *�      ,    ,  .�  *�  R  *�  R  Bh  .�  Bh  .�  *�      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      -    ,  0� �X  S� �X  S� ��  0� ��  0� �X      -    ,  � ��  �� ��  �� ��  � ��  � ��      +    ,  w$  :�  ��  :�  ��  J8  w$  J8  w$  :�      +    ,  �  �  ��  �  ��  #(  �  #(  �  �      +    ,  8� �(  L, �(  L, ��  8� ��  8� �(      +    ,  8� ��  J8 ��  J8 �(  8� �(  8� ��      +    ,  6�  #(  J8  #(  J8  :�  6�  :�  6�  #(      +    ,  8�  :�  HD  :�  HD  J8  8�  J8  8�  :�      +    ,  u0  #(  ��  #(  ��  :�  u0  :�  u0  #(      +    ,  � ��  �� ��  �� �   � �   � ��      0    ,  D\  |  L,  |  L,  L  D\  L  D\  |      0    ,  [�  |  c�  |  c�  L  [�  L  [�  |      0    ,  s<  |  {  |  {  L  s<  L  s<  |      0    ,  ��  |  �|  |  �|  L  ��  L  ��  |      0    ,  �  |  ��  |  ��  L  �  L  �  |      0    ,  {  ,�  ��  ,�  ��  4�  {  4�  {  ,�      0    ,  ,�  |  4�  |  4�  L  ,�  L  ,�  |      0    ,  �� �t  �| �t  �| �D  �� �D  �� �t      0    ,  s< �t  { �t  { �D  s< �D  s< �t      0    ,  [� �t  c� �t  c� �D  [� �D  [� �t      0    ,  D\ �t  L, �t  L, �D  D\ �D  D\ �t      0    ,  ,� �t  4� �t  4� �D  ,� �D  ,� �t      0    ,  | �t  L �t  L �D  | �D  | �t      0    ,  |  |  L  |  L  L  |  L  |  |      0    ,  >� �  FP �  FP ��  >� ��  >� �      0    ,  <�  ,�  D\  ,�  D\  4�  <�  4�  <�  ,�      0    ,  � �t  �� �t  �� �D  � �D  � �t      .    ,  e�  ��  y  ��  y  �P  e�  �P  e�  ��      .    ,  Bh  ��  U�  ��  U�  �P  Bh  �P  Bh  ��      .    ,  ��  ��  �@  ��  �@  �P  ��  �P  ��  ��   	   .      �   0�  g�  0� �   	   .      �   R �  R  �P   	   .      �   ix �  ix  �P   	   .      �   oT  kl  oT  ��   	   .      �   P  kl  P  ��   	   .      �   ��  kl  ��  ��   	   .      � $  �� �  ��  �`  ��  �`  ��  �P      .    ,  ,�  ��  @t  ��  @t  �p  ,�  �p  ,�  ��      /    ,  kl  ��  s<  ��  s<  �t  kl  �t  kl  ��      /    ,  HD  ��  P  ��  P  �t  HD  �t  HD  ��      /    ,  ��  ��  �d  ��  �d  �t  ��  �t  ��  ��      /    ,  2�  ��  :�  ��  :�  ��  2�  ��  2�  ��      1    ,  :� �  J8 �  J8 ��  :� ��  :� �      1    ,  D\  ��  S�  ��  S�  �\  D\  �\  D\  ��      1    ,  g�  ��  w$  ��  w$  �\  g�  �\  g�  ��      1    ,  y  8�  ��  8�  ��  L,  y  L,  y  8�      1    ,  :� ��  HD ��  HD �  :� �  :� ��      1    ,  8�  '  HD  '  HD  8�  8�  8�  8�  '      1    ,  :�  8�  FP  8�  FP  L,  :�  L,  :�  8�      1    ,  w$  '  ��  '  ��  8�  w$  8�  w$  '      1    ,  ��  ��  �L  ��  �L  �\  ��  �\  ��  ��   	   1      �   !4 |  !4  �P   	   1      � $  !4  [�  !4  oT  L  oT  L  ��      1    ,  .�  ��  >�  ��  >�  �|  .�  �|  .�  ��   	   1      �   >�  ��  �4  ��  �4  _�   	   1      �   _�  _�  _�  ��   	   1      � $  �  ��  ��  ��  �� X  �X X              _�  � GND  +  ,1               _� �8 VDD  +  ,1               L  �� Y  +  ,1               oT  �� A1 +  ,1               L,  �� A0 +  ,1               �|  �� A2 +  ,1               _�  � GND               _� �8 VDD               L  �� Y               oT  �� A1              L,  �� A0              �|  �� A2     �  
   � 	   /  
and02     +    <  ,� �  ,� <h  p <h  p p  L p  L �  ,� � +  ,2       0    ,  L L  % L  %   L   L L      0    ,  L .�  % .�  % 6�  L 6�  L .�      1    ,  d d  ) d  ) :t  d :t  d d +  ,1       .    ,  ,�  �  4�  �  4� �  ,� �  ,�  � +  ,3       .    ,  ,� <h  4� <h  4� F,  ,� F,  ,� <h +  ,4       .    ,  ,� �  4� �  4� <h  ,� <h  ,� �      0    ,  <� �  D\ �  D\ |  <� |  <� �      0    ,  <�   D\   D\ &�  <� &�  <�       1    ,  8� �  HD �  HD *�  8� *�  8� � +  ,5       .    ,  L,  �  S�  �  S� �  L, �  L,  � +  ,6       .    ,  L, <h  S� <h  S� F,  L, F,  L, <h +  ,7       .    ,  L, �  S� �  S� <h  L, <h  L, �      0    ,  [� L  c� L  c�   [�   [� L      0    ,  [� .�  c� .�  c� 6�  [� 6�  [� .�      1    ,  W� d  g� d  g� :t  W� :t  W� d +  ,8       .    ,  m`  �  u0  �  u0 �  m` �  m`  � +  ,9       .    ,  m` ,�  u0 ,�  u0 6�  m` 6�  m` ,� +  ,10      .    ,  m` �  u0 �  u0 ,�  m` ,�  m` �      0    ,  }  �  �� �  �� |  }  |  }  �      0    ,  }    ��   �� &�  }  &�  }        1    ,  y �  �� �  �� *�  y *�  y � +  ,11      +    L  �� �  �� ,�  ix ,�  ix <h  p <h  p p  L p  L �  �� �      *    L  �  �`  � D8  �� D8  �� S�     S�      �   �  �   �  �`  �  �` +  ,13      ,    L  �|  �   �| 4�  qH 4�  qH D8  � D8  � 	�  | 	�  |  �   �|  �       +    ,  u0 �  �� �  �� ,�  u0 ,�  u0 � +  ,12      +    ,  ��  ��  u0  ��  u0  �X  ��  �X  ��  �� +  ,2       0    ,  ��  ��  }   ��  }   �|  ��  �|  ��  ��      1    ,  ��  ��  y  ��  y  �d  ��  �d  ��  �� +  ,1       .    ,  u0  {  m`  {  m`  ��  u0  ��  u0  { +  ,3       .    ,  u0  �X  m`  �X  m`  �  u0  �  u0  �X +  ,4       .    ,  u0  ��  m`  ��  m`  �X  u0  �X  u0  ��      0    ,  c�  s<  [�  s<  [�  {  c�  {  c�  s<      0    ,  c�  ��  [�  ��  [�  �|  c�  �|  c�  ��      1    ,  g�  oT  W�  oT  W�  �d  g�  �d  g�  oT +  ,5       .    ,  S�  c�  L,  c�  L,  m`  S�  m`  S�  c� +  ,6       .    ,  S�  �X  L,  �X  L,  �  S�  �  S�  �X +  ,7       .    ,  S�  m`  L,  m`  L,  �X  S�  �X  S�  m`      .    ,  <�  c�  4�  c�  4�  m`  <�  m`  <�  c� +  ,8       .    ,  <�  �X  4�  �X  4�  �  <�  �  <�  �X +  ,9       .    ,  <�  m`  4�  m`  4�  �X  <�  �X  <�  m`      0    ,  ,�  s<  %  s<  %  {  ,�  {  ,�  s<      0    ,  ,�  ��  %  ��  %  �|  ,�  �|  ,�  ��      1    ,  0�  oT  !4  oT  !4  �d  0�  �d  0�  oT +  ,10      +    <  @  m`  @  �X  ��  �X  ��  ��  ix  ��  ix  m`  @  m`      )    <  �  U�  �  ��  �  ��  �  m`  ��  m`  ��  U�  �  U� +  ,12      -    <  p  e�  p  �(  �|  �(  �|  }   qH  }   qH  e�  p  e�      +    ,  4�  m`  @  m`  @  �X  4�  �X  4�  m` +  ,11   
  via  �  B�         Y�  �   
  via  �  B�         ��  �   
  via  �  B�         #(  �      3    ,  ~�  �P  �|  �P  �|  ��  ~�  ��  ~�  �P      3    ,  P  �P  c�  �P  c�  ��  P  ��  P  �P      3    ,  d  �P  ,�  �P  ,�  ��  d  ��  d  �P      1    ,     ��  � ��  � ��     ��     ��      1    ,          �      �  '      '              1    ,     ��  � ��  � ��     ��     ��      1    ,          �      �  '      '                      ��  � Y  +  ,1               Y�  � A1 +  ,1               #(  � A0 +  ,1               Q  � GND  +  ,1               Q �8 VDD  +  ,1       1    ,  L  �D  ,�  �D  ,�  ��  L  ��  L  �D      1    ,  a�  �  qH  �  qH  ��  a�  ��  a�  �   	   1      �   D\  ��  a�  ��   	   1      �   ��  ��  �� |      1    ,  P  �D  _�  �D  _�  ��  P  ��  P  �D   	   1      � $  *�  �d  *�  �  >�  �  >� �      1    ,  Y�  [�  g�  [�  g�  oT  Y�  oT  Y�  [�      1    ,  W�  '  g�  '  g�  [�  W�  [�  W�  '      1    ,  W� M�  g� M�  g� ��  W� ��  W� M�      1    ,  d M�  ) M�  ) ��  d ��  d M�      1    ,  d :t  ' :t  ' M�  d M�  d :t      1    ,  Y� :t  g� :t  g� M�  Y� M�  Y� :t      +    ,  p  �  ��  �  ��  #(  p  #(  p  �      +    ,  p ��  �� ��  �� �   p �   p ��      +    ,  U�  #(  ix  #(  ix  ]�  U�  ]�  U�  #(      +    ,  W�  ]�  ix  ]�  ix  m`  W�  m`  W�  ]�      +    ,  p <h  ) <h  ) L  p L  p <h      +    ,  W� <h  ix <h  ix L  W� L  W� <h      +    ,  p L  *� L  *� ��  p ��  p L      +    ,  U� L  ix L  ix ��  U� ��  U� L      0    ,  c�  |  kl  |  kl  L  c�  L  c�  |      0    ,  {  |  ��  |  ��  L  {  L  {  |      0    ,  L,  |  S�  |  S�  L  L,  L  L,  |      0    ,  { �t  �� �t  �� �D  { �D  { �t      0    ,  4�  |  <�  |  <�  L  4�  L  4�  |      0    ,  L  |  %  |  %  L  L  L  L  |      0    ,  4� �t  <� �t  <� �D  4� �D  4� �t      0    ,  L, �t  S� �t  S� �D  L, �D  L, �t      0    ,  c� �t  kl �t  kl �D  c� �D  c� �t      0    ,  L �t  % �t  % �D  L �D  L �t      0    ,  [�  P  c�  P  c�  W�  [�  W�  [�  P      0    ,  [�  8�  c�  8�  c�  @t  [�  @t  [�  8�      0    ,  [� iT  c� iT  c� q$  [� q$  [� iT      0    ,  [� ��  c� ��  c� ��  [� ��  [� ��      0    ,  [� �4  c� �4  c� �  [� �  [� �4      0    ,  L ��  % ��  % ��  L ��  L ��      0    ,  L iT  % iT  % q$  L q$  L iT      0    ,  [� Q�  c� Q�  c� Y�  [� Y�  [� Q�      0    ,  L Q�  % Q�  % Y�  L Y�  L Q�      0    ,  L �4  % �4  % �  L �  L �4      -    ,  � ��  �� ��  �� ��  � ��  � ��      -    ,  N  D8  qH D8  qH ��  N  ��  N  D8      -    ,  � D8  2� D8  2� ��  � ��  � D8      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      ,    ,  N   *�  qH  *�  qH  e�  N   e�  N   *�      )    ,          �      �  ��      ��              *    ,      �`  �  �`  � ��     ��      �`      .    ,  _�  �(  s<  �(  s<  ��  _�  ��  _�  �(   	   .      �   P  �  P  �   	   .      �   0�  �  0�  �  <�  �   	   .      �   qH  �  qH  �      .    ,  N   �P  a�  �P  a�  ��  N   ��  N   �P      .    ,  X  �P  .�  �P  .�  ��  X  ��  X  �P      /    ,  e�  �  m`  �  m`  ��  e�  ��  e�  �      /    ,  S�  �,  [�  �,  [�  ��  S�  ��  S�  �,      /    ,  !4  �,  )  �,  )  ��  !4  ��  !4  �,      �    ,          �      � ��     ��                      Q  � GND               Q �8 VDD               ��  � Y               Y�  � A1              #(  � A0     �    4 � 	   / 8 dffr    0    , �\ :t �� :t �� BD �\ BD �\ :t      0    , �\ Q� �� Q� �� Y� �\ Y� �\ Q�      0    , �\ iT �� iT �� q$ �\ q$ �\ iT      1    , �D 6� �� 6� �� u �D u �D 6� +  ,1       .    , �� *� �� *� �� 4� �� 4� �� *� +  ,3       .    , �� �� �� �� �� �L �� �L �� �� +  ,4       .    , �� 4� �� 4� �� �� �� �� �� 4�      0    , � M� �L M� �L U� � U� � M�      0    , � el �L el �L m< � m< � el      0    , � |� �L |� �L �� � �� � |�      1    , � J �d J �d �� � �� � J +  ,5       .    , �| *� ~� *� ~� 4� �| 4� �| *� +  ,6       .    , �| �� ~� �� ~� �L �| �L �| �� +  ,7       .    , �| 4� ~� 4� ~� �� �| �� �| 4�      0    , v� :t o :t o BD v� BD v� :t      0    , v� Q� o Q� o Y� v� Y� v� Q�      0    , v� iT o iT o q$ v� q$ v� iT      1    , z� 6� k$ 6� k$ u z� u z� 6� +  ,8       +    L i0 4� i0 w  o w  o �� �\ �� �\ w  �8 w  �8 4� i0 4�      *    L Q� ( Q� �p W� �p W� �� �� �� �� �p Ҩ �p Ҩ ( Q� ( +  ,10      ,    L a` ,� a` ~� g< ~� g< �X �, �X �, ~� � ~� � ,� a` ,�      +    < i0 4� i0 w  o w  o �� ~� �� ~� 4� i0 4� +  ,9       +    < �� 4� �� �� �\ �� �\ w  �8 w  �8 4� �� 4� +  ,2       +    , p J  �� J  �� u p u p J +  ,2       0    , � O� � O� � W� � W� � O�      0    , � g` � g` � o0 � o0 � g`      1    , | L  �� L  �� s | s | L +  ,1       .    ,  �� @P  �$ @P  �$ J  �� J  �� @P +  ,3       .    ,  �� u  �$ u  �$ ~�  �� ~�  �� u +  ,4       .    ,  �� J  �$ J  �$ u  �� u  �� J      0    ,  �T O�  � O�  � W�  �T W�  �T O�      0    ,  �T g`  � g`  � o0  �T o0  �T g`      1    ,  �< L  �� L  �� s  �< s  �< L +  ,5       +    , p J  ި J  ި u p u p J      *    , (� 2�  �8 2�  �8 �| (� �| (� 2� +  ,7       ,    , @ BD  �� BD  �� |� @ |� @ BD      +    ,  �$ J  ި J  ި u  �$ u  �$ J +  ,6       0    ,  L   %   % &�  L &�  L       0    ,  L 6�  % 6�  % >\  L >\  L 6�      0    ,  L M�  % M�  % U�  L U�  L M�      0    ,  L el  % el  % m<  L m<  L el      0    ,  L |�  % |�  % ��  L ��  L |�      1    ,  d 4  ) 4  ) ��  d ��  d 4 +  ,1       .    ,  ,� �  4� �  4� �  ,� �  ,� � +  ,3       .    ,  ,� ��  4� ��  4� �L  ,� �L  ,� �� +  ,4       .    ,  ,� �  4� �  4� ��  ,� ��  ,� �      .    ,  D\ �  L, �  L, �  D\ �  D\ � +  ,5       .    ,  D\ ��  L, ��  L, �L  D\ �L  D\ �� +  ,6       .    ,  D\ �  L, �  L, ��  D\ ��  D\ �      0    ,  S� d  [� d  [� 4  S� 4  S� d      0    ,  S� *�  [� *�  [� 2�  S� 2�  S� *�      0    ,  S� BD  [� BD  [� J  S� J  S� BD      0    ,  S� Y�  [� Y�  [� a�  S� a�  S� Y�      0    ,  S� q$  [� q$  [� x�  S� x�  S� q$      1    ,  P |  _� |  _� |�  P |�  P | +  ,7       .    ,  e� W�  m` W�  m` a�  e� a�  e� W� +  ,8       .    ,  e� u  m` u  m` ~�  e� ~�  e� u +  ,9       .    ,  e� a�  m` a�  m` u  e� u  e� a�      .    ,  }  W�  �� W�  �� a�  }  a�  }  W� +  ,10      .    ,  }  u  �� u  �� ~�  }  ~�  }  u +  ,11      .    ,  }  a�  �� a�  �� u  }  u  }  a�      0    ,  �� O�  �d O�  �d W�  �� W�  �� O�      0    ,  �� g`  �d g`  �d o0  �� o0  �� g`      1    ,  �� L  �L L  �L s  �� s  �� L +  ,12      .    ,  �4 0�  � 0�  � :t  �4 :t  �4 0� +  ,13      .    ,  �4 u  � u  � ~�  �4 ~�  �4 u +  ,14      .    ,  �4 :t  � :t  � u  �4 u  �4 :t      .    ,  �� 0�  �t 0�  �t :t  �� :t  �� 0� +  ,15      .    ,  �� u  �t u  �t ~�  �� ~�  �� u +  ,16      .    ,  �� :t  �t :t  �t u  �� u  �� :t      0    ,  �D @P  � @P  � H   �D H   �D @P      0    ,  �D W�  � W�  � _�  �D _�  �D W�      1    ,  �\ <h  �� <h  �� cx  �\ cx  �\ <h +  ,17      +    �  a� �  a� a�  �� a�  �� J  �� J  �� :t  �� :t  �� el  � el  � u  a� u  a� ~�  [� ~�  [� ��  p ��  p @  L @  L �  a� �      *    |  y  �  y #  �` #  �` |�  � |�  � �|  y �|  y �@  s< �@  s< ��     ��     �  � �  �  �  y  � +  ,19      ,    �  ix �  ix Y�  �� Y�  �� BD  �� BD  �� 2�  �� 2�  �� m<  �� m<  �� |�  ix |�  ix ��  c� ��  c� �X  � �X  � p  | p  | �  ix �      +    <  �� :t  �� el  � el  � u  �t u  �t :t  �� :t +  ,18      +    <  ,� �  ,� ��  p ��  p @  L @  L �  ,� � +  ,2       +    , (  �� 2�  �� 2�  �� (  �� (  �� +  ,2       0    , #  �� *�  �� *�  �� #  �� #  ��      0    , #  �4 *�  �4 *�  � #  � #  �4      1    ,   �� .�  �� .�  ��   ��   �� +  ,1       .    , 2�  w$ :t  w$ :t  �� 2�  �� 2�  w$ +  ,3       .    , 2�  �� :t  �� :t  �� 2�  �� 2�  �� +  ,4       .    , 2�  �� :t  �� :t  �� 2�  �� 2�  ��      0    , BD  �� J  �� J  �� BD  �� BD  ��      0    , BD  �4 J  �4 J  � BD  � BD  �4      1    , >\  �� M�  �� M�  �� >\  �� >\  �� +  ,5       .    , Q�  w$ Y�  w$ Y�  �� Q�  �� Q�  w$ +  ,6       .    , Q�  �� Y�  �� Y�  �� Q�  �� Q�  �� +  ,7       .    , Q�  �� Y�  �� Y�  �� Q�  �� Q�  ��      0    , a�  �� iT  �� iT  �� a�  �� a�  ��      0    , a�  �4 iT  �4 iT  � a�  � a�  �4      1    , ]�  �� m<  �� m<  �� ]�  �� ]�  �� +  ,8       +    , (  �� o0  �� o0  �� (  �� (  ��      )    , �  ix ��  ix ��  �P �  �P �  ix +  ,10      -    , X  y w   y w   �� X  �� X  y      +    , Y�  �� o0  �� o0  �� Y�  �� Y�  �� +  ,9       0    ,  �  ��  �H  ��  �H  ��  �  ��  �  ��      1    ,  �   ��  �`  ��  �`  �|  �   �|  �   �� +  ,1       .    ,  �x  w$  ި  w$  ި  ��  �x  ��  �x  w$ +  ,3       .    ,  �x  �p  ި  �p  ި  �4  �x  �4  �x  �p +  ,4       .    ,  �x  ��  ި  ��  ި  �p  �x  �p  �x  ��      0    ,  ��  oT  �  oT  �  w$  ��  w$  ��  oT      0    ,  ��  ��  �  ��  �  ��  ��  ��  ��  ��      1    ,  ��  kl  �,  kl  �,  �|  ��  �|  ��  kl +  ,5       .    ,  �D  _�  �t  _�  �t  ix  �D  ix  �D  _� +  ,6       .    ,  �D  �p  �t  �p  �t  �4  �D  �4  �D  �p +  ,7       .    ,  �D  ix  �t  ix  �t  �p  �D  �p  �D  ix      0    ,  ��  oT  ��  oT  ��  w$  ��  w$  ��  oT      0    ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��      1    ,  ��  kl  ��  kl  ��  �|  ��  �|  ��  kl +  ,8       .    ,  �  _�  �4  _�  �4  ix  �  ix  �  _� +  ,9       .    ,  �  �p  �4  �p  �4  �4  �  �4  �  �p +  ,10      .    ,  �  ix  �4  ix  �4  �p  �  �p  �  ix      0    ,  �d  oT  ��  oT  ��  w$  �d  w$  �d  oT      0    ,  �d  ��  ��  ��  ��  ��  �d  ��  �d  ��      1    ,  �L  kl  ��  kl  ��  �|  �L  �|  �L  kl +  ,11      .    ,  ��  w$  }   w$  }   ��  ��  ��  ��  w$ +  ,12      .    ,  ��  �p  }   �p  }   �4  ��  �4  ��  �p +  ,13      .    ,  ��  ��  }   ��  }   �p  ��  �p  ��  ��      .    ,  m`  w$  e�  w$  e�  ��  m`  ��  m`  w$ +  ,14      .    ,  m`  �p  e�  �p  e�  �4  m`  �4  m`  �p +  ,15      .    ,  m`  ��  e�  ��  e�  �p  m`  �p  m`  ��      0    ,  [�  W�  S�  W�  S�  _�  [�  _�  [�  W�      0    ,  [�  oT  S�  oT  S�  w$  [�  w$  [�  oT      0    ,  [�  ��  S�  ��  S�  ��  [�  ��  [�  ��      1    ,  _�  S�  P  S�  P  �|  _�  �|  _�  S� +  ,16      .    ,  L,  HD  D\  HD  D\  R  L,  R  L,  HD +  ,17      .    ,  L,  �p  D\  �p  D\  �4  L,  �4  L,  �p +  ,18      .    ,  L,  R  D\  R  D\  �p  L,  �p  L,  R      .    ,  4�  HD  ,�  HD  ,�  R  4�  R  4�  HD +  ,19      .    ,  4�  �p  ,�  �p  ,�  �4  4�  �4  4�  �p +  ,20      .    ,  4�  R  ,�  R  ,�  �p  4�  �p  4�  R      0    ,  %  W�  L  W�  L  _�  %  _�  %  W�      0    ,  %  oT  L  oT  L  w$  %  w$  %  oT      0    ,  %  ��  L  ��  L  ��  %  ��  %  ��      1    ,  )  S�  d  S�  d  �|  )  �|  )  S� +  ,21      +    \  p  R  p  �p  ��  �p  ��  ��  ��  ��  ��  ix  ��  ix  ��  ��  a�  ��  a�  R  p  R      )    L      :�      �� d  �� d  ix  �0  ix  �0  R  y  R  y  :�      :� +  ,23      -    \  �  J8  �  �@ �  �@ �  y  �  y  �  a�  ��  a�  ��  y  ix  y  ix  J8  �  J8      +    ,  ,�  R  p  R  p  �p  ,�  �p  ,�  R +  ,22      +    ,  ��  ��  �x  ��  �x  �p  ��  �p  ��  �� +  ,2       +    , (� _� >8 _� >8 �� (� �� (� _� +  ,2       0    , .� el 6h el 6h m< .� m< .� el      0    , .� |� 6h |� 6h �� .� �� .� |�      1    , *� a� :P a� :P �� *� �� *� a� +  ,1       .    , >8 U� F U� F _� >8 _� >8 U� +  ,3       .    , >8 �� F �� F �L >8 �L >8 �� +  ,4       .    , >8 _� F _� F �� >8 �� >8 _�      0    , M� el U� el U� m< M� m< M� el      0    , M� |� U� |� U� �� M� �� M� |�      1    , I� a� Y� a� Y� �� I� �� I� a� +  ,5       +    , (� _� [� _� [� �� (� �� (� _�      *    , L H  r� H  r� �� L �� L H  +  ,7       ,    ,  � W� cT W� cT �X  � �X  � W�      +    , F _� [� _� [� �� F �� F _� +  ,6       0    , .� d &� d &� 4 .� 4 .� d      1    , 2� | "� | "�  2�  2� | +  ,1       .    , � � ( � ( � � � � � +  ,3       .    , � ! ( ! ( *� � *� � ! +  ,4       .    , � � ( � ( ! � ! � �      .    , � � �� � �� � � � � � +  ,5       .    , � ! �� ! �� *� � *� � ! +  ,6       .    , � � �� � �� ! � ! � �      0    , ��  �$  �$ &� �� &� ��       0    , �� 6� �$ 6� �$ >\ �� >\ �� 6�      0    , �� M� �$ M� �$ U� �� U� �� M�      0    , �� el �$ el �$ m< �� m< �� el      0    , �� |� �$ |� �$ �� �� �� �� |�      1    , �� 4 �< 4 �< �� �� �� �� 4 +  ,7       .    , �T � ބ � ބ � �T � �T � +  ,8       .    , �T �� ބ �� ބ �L �T �L �T �� +  ,9       .    , �T � ބ � ބ �� �T �� �T �      .    , �� � � � � � �� � �� � +  ,10      .    , �� �� � �� � �L �� �L �� �� +  ,11      .    , �� � � � � �� �� �� �� �      0    , �D  �t  �t &� �D &� �D       0    , �D 6� �t 6� �t >\ �D >\ �D 6�      0    , �D M� �t M� �t U� �D U� �D M�      0    , �D el �t el �t m< �D m< �D el      0    , �D |� �t |� �t �� �D �� �D |�      1    , �, 4 �� 4 �� �� �, �� �, 4 +  ,12      .    , �� � �� � �� � �� � �� � +  ,13      .    , �� ! �� ! �� *� �� *� �� ! +  ,14      .    , �� � �� � �� ! �� ! �� �      0    , � d �@ d �@ 4 � 4 � d      1    , �� | �X | �X  ��  �� | +  ,15      +    L �d � �d ! �� ! �� �� �� �� �� ! 4t ! 4t � �d �      *    L x�  � x� 8� �( 8� �( �� @ �� @ 8� K� 8� K�  � x�  � +  ,17      ,    L �� � �� (� �� (� �� �X � �X � (� <D (� <D � �� �      +    , �� � �d � �d ! �� ! �� � +  ,16      +    , 4t � � � � ! 4t ! 4t � +  ,2       0    , iT &� a� &� a� .� iT .� iT &�      0    , iT >\ a� >\ a� F, iT F, iT >\      0    , iT U� a� U� a� ]� iT ]� iT U�      1    , m< # ]� # ]� a� m< a� m< # +  ,1       .    , Y� L Q� L Q� ! Y� ! Y� L +  ,3       .    , Y� w  Q� w  Q� �� Y� �� Y� w  +  ,4       .    , Y� ! Q� ! Q� w  Y� w  Y� !      0    , J :t BD :t BD BD J BD J :t      0    , J Q� BD Q� BD Y� J Y� J Q�      0    , J iT BD iT BD q$ J q$ J iT      1    , M� 6� >\ 6� >\ u M� u M� 6� +  ,5       .    , :t L 2� L 2� ! :t ! :t L +  ,6       .    , :t w  2� w  2� �� :t �� :t w  +  ,7       .    , :t ! 2� ! 2� w  :t w  :t !      0    , *� &� # &� # .� *� .� *� &�      0    , *� >\ # >\ # F, *� F, *� >\      0    , *� U� # U� # ]� *� ]� *� U�      1    , .� #  #  a� .� a� .� # +  ,8       +    L ( ! ( cx # cx # w  iT w  iT cx o0 cx o0 ! ( !      *    L � 	� � z� � z� � �p �� �p �� z� �� z� �� 	� � 	� +  ,10      ,    L X @ X kH 4 kH 4 ~� q$ ~� q$ kH w  kH w  @ X @      +    < ( ! ( cx # cx # w  2� w  2� ! ( ! +  ,9       +    < Y� ! Y� w  iT w  iT cx o0 cx o0 ! Y� ! +  ,2       0    , U�  ix M�  ix M�  qH U�  qH U�  ix      1    , Y�  e� I�  e� I�  u0 Y�  u0 Y�  e� +  ,1       .    , F  Y� >8  Y� >8  c� F  c� F  Y� +  ,3       .    , F  w$ >8  w$ >8  �� F  �� F  w$ +  ,4       .    , F  c� >8  c� >8  w$ F  w$ F  c�      0    , 6h  ix .�  ix .�  qH 6h  qH 6h  ix      1    , :P  e� *�  e� *�  u0 :P  u0 :P  e� +  ,5       .    , &�  Y� �  Y� �  c� &�  c� &�  Y� +  ,6       .    , &�  w$ �  w$ �  �� &�  �� &�  w$ +  ,7       .    , &�  c� �  c� �  w$ &�  w$ &�  c�      0    , (  ix X  ix X  qH (  qH (  ix      1    ,   e� p  e� p  u0   u0   e� +  ,8       .    , �  Y� ��  Y� ��  c� �  c� �  Y� +  ,9       .    , �  w$ ��  w$ ��  �� �  �� �  w$ +  ,10      .    , �  c� ��  c� ��  w$ �  w$ �  c�      0    , ��  ix �$  ix �$  qH ��  qH ��  ix      0    , ��  �� �$  �� �$  �� ��  �� ��  ��      0    , ��  �X �$  �X �$  �( ��  �( ��  �X      1    , ��  e� �<  e� �<  � ��  � ��  e� +  ,11      .    , �T  Y� ބ  Y� ބ  c� �T  c� �T  Y� +  ,12      .    , �T  � ބ  � ބ  �� �T  �� �T  � +  ,13      .    , �T  c� ބ  c� ބ  � �T  � �T  c�      .    , ��  Y� �  Y� �  c� ��  c� ��  Y� +  ,14      .    , ��  � �  � �  �� ��  �� ��  � +  ,15      .    , ��  c� �  c� �  � ��  � ��  c�      0    , �D  ix �t  ix �t  qH �D  qH �D  ix      0    , �D  �� �t  �� �t  �� �D  �� �D  ��      0    , �D  �X �t  �X �t  �( �D  �( �D  �X      1    , �,  e� ��  e� ��  � �,  � �,  e� +  ,16      .    , ��  �� ��  �� ��  �| ��  �| ��  �� +  ,17      .    , ��  � ��  � ��  �� ��  �� ��  � +  ,18      .    , ��  �| ��  �| ��  � ��  � ��  �|      0    , �  �X �@  �X �@  �( �  �( �  �X      1    , ��  �p �X  �p �X  � ��  � ��  �p +  ,19      +    L ��  c� ��  �| �d  �| �d  � ��  � ��  w$ [�  w$ [�  c� ��  c�      )    L �(  L, �(  { x�  { x�  �t @  �t @  �� r�  �� r�  L, �(  L, +  ,21      -    L ��  [� ��  �� ��  �� ��  �� �  �� �  ~� cT  ~� cT  [� ��  [�      +    , ��  �| �d  �| �d  � ��  � ��  �| +  ,20      +    , [�  c� F  c� F  w$ [�  w$ [�  c� +  ,2       +    , �8  J8 ��  J8 ��  u0 �8  u0 �8  J8 +  ,2       0    , �\  P ��  P ��  W� �\  W� �\  P      0    , �\  g� ��  g� ��  oT �\  oT �\  g�      1    , �D  L, ��  L, ��  s< �D  s< �D  L, +  ,1       .    , ��  @t ��  @t ��  J8 ��  J8 ��  @t +  ,3       .    , ��  u0 ��  u0 ��  ~� ��  ~� ��  u0 +  ,4       .    , ��  J8 ��  J8 ��  u0 ��  u0 ��  J8      0    , �  P �L  P �L  W� �  W� �  P      0    , �  g� �L  g� �L  oT �  oT �  g�      1    , �  L, �d  L, �d  s< �  s< �  L, +  ,5       .    , �|  @t ~�  @t ~�  J8 �|  J8 �|  @t +  ,6       .    , �|  u0 ~�  u0 ~�  ~� �|  ~� �|  u0 +  ,7       .    , �|  J8 ~�  J8 ~�  u0 �|  u0 �|  J8      0    , v�  P o  P o  W� v�  W� v�  P      0    , v�  g� o  g� o  oT v�  oT v�  g�      1    , z�  L, k$  L, k$  s< z�  s< z�  L, +  ,8       +    , �8  J8 i0  J8 i0  u0 �8  u0 �8  J8      )    , Ҩ  2� Q�  2� Q�  �� Ҩ  �� Ҩ  2� +  ,10      -    , �  Bh a`  Bh a`  }  �  }  �  Bh      +    , ~�  J8 i0  J8 i0  u0 ~�  u0 ~�  J8 +  ,9    
  via  �  B�        �\  �   
  via  �  B�        >\  �   
  via  �  B�         �  �   
  via  �  B�         Bh  �   
  via  �  B�        q   �      3    ,  �D  �P  ��  �P  ��  ��  �D  ��  �D  �P      3    ,  8�  �P  L,  �P  L,  ��  8�  ��  8�  �P      3    , 4�  �P H   �P H   �� 4�  �� 4�  �P      3    , ��  �P �   �P �   �� ��  �� ��  �P      3    , g<  �P z�  �P z�  �� g<  �� g<  �P      1    ,     �� Ҩ �� Ҩ ��     ��     ��      1    ,         Ҩ     Ҩ  '      '              �    ,         Ҩ     Ҩ ��     ��                     n6  � GND  +  ,1       /    ,  �,  �,  ��  �,  ��  ��  �,  ��  �,  �,      /    , �  �� �  �� �  �� �  �� �  ��      /    , �x  ܴ �H  ܴ �H  � �x  � �x  ܴ      /    ,  >�  �,  FP  �,  FP  ��  >�  ��  >�  �,      /    , #  6� *�  6� *�  >� #  >� #  6�      /    , ��  ܴ ��  ܴ ��  � ��  � ��  ܴ      /    , a�  FP iT  FP iT  N  a�  N  a�  FP      /    ,  _�  �x  g�  �x  g�  �H  _�  �H  _�  �x      /    ,  ��  �,  �X  �,  �X  ��  ��  ��  ��  �,      /    ,  ��  D\  ��  D\  ��  L,  ��  L,  ��  D\      /    ,  '  �  .�  �  .�  ��  '  ��  '  �      /    , L  �0 S�  �0 S�  �  L  �  L  �0      /    , 8�  �, @P  �, @P  �� 8�  �� 8�  �,      /    , �  ܴ 	|  ܴ 	|  � �  � �  ܴ   	   .      �   ix  w$  ix  HD  ��  HD      .    , ��  �� X  �� X  �` ��  �` ��  ��   	   .      �  Y�  �� ��  ��   	   .      �  ��  �� ��  �`      .    , ڜ  �� �$  �� �$  �` ڜ  �` ڜ  ��      .    , [�  @t o0  @t o0  S� [�  S� [�  @t   	   .      � , �l  Y� �l  Bh ��  Bh ��  D\ o0  D\   	   .      � <  �t  a�  �`  a�  �`  S� F,  S� F,  .� "�  .� "�  0�      .    , ��  �� �\  �� �\  �` ��  �` ��  ��      .    ,  ��  �� d  �� d  �p  ��  �p  ��  ��      .    , (  0� 0�  0� 0�  D\ (  D\ (  0�      .    ,  8�  �P  L,  �P  L,  ��  8�  ��  8�  �P   	   .      �   0�  HD  0�  .� 0�  .�   	   .      � $  ��  �4  ��  ��  ix  ��  ix  ��      .    ,  Y�  ��  m`  ��  m`  �$  Y�  �$  Y�  ��      .    ,  ��  �P  �4  �P  �4  ��  ��  ��  ��  �P   	   .      � $  �  �4  �  �  �`  �  �`  �      .    , F,  �T Y�  �T Y�  �� F,  �� F,  �T      .    ,  �P  �P  ��  �P  ��  ��  �P  ��  �P  �P      .    ,  ��  >�  ��  >�  ��  R  ��  R  ��  >�   	   .      � 4 |  �� |  g� ��  g� ��  U� ��  U� ��  Y�      .    , 2�  �P F,  �P F,  �� 2�  �� 2�  �P   	   .      �  "�  0� "�  Y�      ,    ,  �  � �  � �  *�  �  *�  �  �      ,    ,  �  *�  0�  *�  0�  J8  �  J8  �  *�      ,    , �l  *� �  *� �  [� �l  [� �l  *�      ,    , "�  *� F  *� F  [� "�  [� "�  *�      ,    , ��  *� ��  *� ��  Bh ��  Bh ��  *�      0    ,  X  |  #(  |  #(  L  X  L  X  |      0    , |�  | ��  | ��  L |�  L |�  |      0    , 0�  D\ 8\  D\ 8\  L, 0�  L, 0�  D\      0    , ��  | �h  | �h  L ��  L ��  |      0    , 0�  ,� 8\  ,� 8\  4� 0�  4� 0�  ,�      0    , �  HD ��  HD ��  P �  P �  HD      0    ,  2�  |  :�  |  :�  L  2�  L  2�  |      0    ,  X  0�  #(  0�  #(  8�  X  8�  X  0�      0    , �(  | ��  | ��  L �(  L �(  |      0    , eH  | m  | m  L eH  L eH  |      0    , M�  | U�  | U�  L M�  L M�  |      0    , 6h  | >8  | >8  L 6h  L 6h  |      0    , �  | &�  | &�  L �  L �  |      0    , �  | X  | X  L �  L �  |      0    , �  | ��  | ��  L �  L �  |      0    , ب  | �x  | �x  L ب  L ب  |      0    , �8  | �  | �  L �8  L �8  |      0    , ��  | ��  | ��  L ��  L ��  |      0    , �X  | �(  | �(  L �X  L �X  |      0    , z�  | ��  | ��  L z�  L z�  |      0    , cx  | kH  | kH  L cx  L cx  |      0    , L  | S�  | S�  L L  L L  |      0    , 4�  | <h  | <h  L 4�  L 4�  |      0    , (  | $�  | $�  L (  L (  |      0    , �  | �  | �  L �  L �  |      0    ,  �H  |  �  |  �  L  �H  L  �H  |      0    ,  ��  |  ި  |  ި  L  ��  L  ��  |      0    ,  �h  |  �8  |  �8  L  �h  L  �h  |      0    ,  ��  |  ��  |  ��  L  ��  L  ��  |      0    ,  ��  |  �X  |  �X  L  ��  L  ��  |      0    ,  y  |  ��  |  ��  L  y  L  y  |      0    ,  a�  |  ix  |  ix  L  a�  L  a�  |      0    ,  J8  |  R  |  R  L  J8  L  J8  |      0    , �L  ,� �  ,� �  4� �L  4� �L  ,�      +    ,  p  D\  )  D\  )  R  p  R  p  D\      +    ,  |  #(  )  #(  )  D\  |  D\  |  #(      +    ,  |  � �D  � �D  #(  |  #(  |  �      +    , *�  #( >8  #( >8  S� *�  S� *�  #(      +    , �p  #( ��  #( ��  :� �p  :� �p  #(      +    , *�  S� :P  S� :P  c� *�  c� *�  S�      +    , �<  U� ��  U� ��  c� �<  c� �<  U�      +    , �<  Bh ��  Bh ��  U� �<  U� �<  Bh      +    , �d  :� �  :� �  J8 �d  J8 �d  :�   	   1      �  �  D\ �  '      1    , ��  �� d  �� d  �l ��  �l ��  ��      1    , ܐ  �� �0  �� �0  �l ܐ  �l ܐ  ��      1    , �  �� p  �� p  �| �  �| �  ��      1    ,  ��  @t  ��  @t  ��  P  ��  P  ��  @t      1    , �d  ' �  ' �  8� �d  8� �d  '      1    , ]�  Bh m<  Bh m<  R ]�  R ]�  Bh   	   1      � $ �  � �  �� L  �� L  u0   	   1      �  K�  �� d  ��      1    , ,�  R 8\  R 8\  e� ,�  e� ,�  R      1    , �0  S� ��  S� ��  e� �0  e� �0  S�      1    , ��  �� �h  �� �h  �l ��  �l ��  ��   	   1      �  F,  �� F,  '      1    ,   2� .�  2� .�  Bh   Bh   2�   	   1      �  ܐ  �� �h  ��   	   1      �   �   �� �  ��   	   1      �  &�  �� &�  Bh      1    ,  p  '  '  '  '  Bh  p  Bh  p  '   	   1      �  el  R el  ��   	   1      �  H   � (�  �   	   1      �   �|  kl  �|  '   	   1      �   ��  kl  ��  '      1    , ,�  ' <D  ' <D  R ,�  R ,�  '      1    ,  [�  �  kl  �  kl  �0  [�  �0  [�  �      1    ,  ��  �D  �@  �D  �@  ��  ��  ��  ��  �D      1    ,  d  Bh  '  Bh  '  S�  d  S�  d  Bh   	   1      �   [�  �T  ,�  �T  ,�  �$      1    ,  :�  �D  J8  �D  J8  ��  :�  ��  :�  �D      1    ,  �D  �D  ��  �D  ��  ��  �D  ��  �D  �D      1    , H   �H W�  �H W�  �� H   �� H   �H      1    , �0  D\ ��  D\ ��  S� �0  S� �0  D\      1    , 4�  �D D8  �D D8  �� 4�  �� 4�  �D   	   1      �   ��  kl  ��  P      1    , �X  8� �  8� �  L, �X  L, �X  8�              �  � R  +  ,1               Bh  � D  +  ,1              >\  � CLK  +  ,1              �\  � Q  +  ,1              q   � QB +  ,1       )    ,         Ҩ     Ҩ  �P      �P                     n6 �8 VDD  +  ,1       -    ,  � �X  0� �X  0� ��  � ��  � �X      -    ,  � �� � �� � ��  � ��  � ��      -    , 4� ~� W� ~� W� �� 4� �� 4� ~�      -    , � W�  � W�  � �X � �X � W�      -    , � �X B  �X B  �� � �� � �X      -    , �� �X �� �X �� �� �� �� �� �X      0    , �� �t �h �t �h �D �� �D �� �t      0    ,  X �t  #( �t  #( �D  X �D  X �t      0    ,  2� �t  :� �t  :� �D  2� �D  2� �t      0    , BD �| J �| J �L BD �L BD �|      0    , 	| el L el L m< 	| m< 	| el      0    ,  X �  #( �  #( ��  X ��  X �      0    , �( �t �� �t �� �D �( �D �( �t      0    , |� �t �� �t �� �D |� �D |� �t      0    , eH �t m �t m �D eH �D eH �t      0    , M� �t U� �t U� �D M� �D M� �t      0    , 6h �t >8 �t >8 �D 6h �D 6h �t      0    , � �t &� �t &� �D � �D � �t      0    , � �t X �t X �D � �D � �t      0    , � �t �� �t �� �D � �D � �t      0    , ب �t �x �t �x �D ب �D ب �t      0    , �8 �t � �t � �D �8 �D �8 �t      0    , �� �t �� �t �� �D �� �D �� �t      0    , �X �t �( �t �( �D �X �D �X �t      0    , z� �t �� �t �� �D z� �D z� �t      0    , cx �t kH �t kH �D cx �D cx �t      0    , L �t S� �t S� �D L �D L �t      0    , 4� �t <h �t <h �D 4� �D 4� �t      0    , ( �t $� �t $� �D ( �D ( �t      0    , � �t � �t � �D � �D � �t      0    ,  �H �t  � �t  � �D  �H �D  �H �t      0    ,  �� �t  ި �t  ި �D  �� �D  �� �t      0    ,  �h �t  �8 �t  �8 �D  �h �D  �h �t      0    ,  �� �t  �� �t  �� �D  �� �D  �� �t      0    ,  �� �t  �X �t  �X �D  �� �D  �� �t      0    ,  y �t  �� �t  �� �D  y �D  y �t      0    ,  a� �t  ix �t  ix �D  a� �D  a� �t      0    ,  J8 �t  R �t  R �D  J8 �D  J8 �t      0    , 	| |� L |� L �� 	| �� 	| |�      0    , ,� � 4t � 4t �� ,� �� ,� �      0    , �L � � � � �� �L �� �L �      +    , �� _� ( _� ( �� �� �� �� _�      +    ,  | �� �D �� �D �   | �   | ��      +    , >\ w  M� w  M� �� >\ �� >\ w       +    , &� �( :P �( :P �� &� �� &� �(      +    , <h �� O� �� O� �( <h �( <h ��      +    , �p �( �� �( �� �� �p �� �p �(      +    ,  | �(  ) �(  ) ��  | ��  | �(      +    ,  p ��  ) ��  ) �(  p �(  p ��      +    , (� �� :P �� :P �( (� �( (� ��      +    , �d �� � �� � �( �d �( �d ��      /    ,  ��  ��  �l  ��  �l �  �� �  ��  ��      /    , �� �@ �� �@ �� � �� � �� �@      /    , �� M� �� M� �� U� �� U� �� M�      /    , _� �@ g` �@ g` � _� � _� �@      /    ,  qH 4�  y 4�  y <h  qH <h  qH 4�      /    , @ �� ! �� ! �d @ �d @ ��      /    , � � �� � �� | � | � �   	   .      �  6� L 6�  ��      .    , �4 � �� � �� X �4 X �4 �   	   .      �  ��  ~� �� *�   	   .      �  �� � ��  ��   	   .      �   ix W�  ix .�   	   .      �  �� *� ��  }       .    , z� H  �p H  �p [� z� [� z� H    	   .      �  � � �  ��   	   .      �  "�  �� "� � ( �   	   .      � $  �` 	�  �` 8�  � 8�  � @P   	   .      � , >8 D8 � D8 � �� �� �� �� ��   	   .      �  �� *� �� L �p L   	   .      �  d �X  �� �X  �� ~�      .    , Y� �d m< �d m< �� Y� �� Y� �d   	   .      �   HD �  HD  �4      .    , �� �d �h �d �h �� �� �� �� �d      .    ,  kl .�  ~� .�  ~� BD  kl BD  kl .�      .    ,  !4  �0  4�  �0  4� �  !4 �  !4  �0   	   .      �  B  U� B   ��   	   .      �  U�  �� U� L   	   .      �   �  �4  � 0�   	   .      � $  �� 0�  �� &�  �\ &�  �\  �4   	   .      �   0� �L  0� �� m< ��   	   .      �  �l � �l  �`      .    , d �� &� �� &� �@ d �@ d ��      .    ,  ��  �  �H  �  �H 	�  �� 	�  ��  �   	   .      �  ~� &� F &�   	   1      � $ (� | (� � � � � |      1    ,  ܴ  �  �T  �  �T �  ܴ �  ܴ  �      1    , �� a� 4 a� 4 �� �� �� �� a�   	   1      �   �D  ��  ��  ��  ��  �|   	   1      �  �( � t� �   	   1      �   �| s  �| ��      1    , @P u L u L �� @P �� @P u   	   1      �  �� �X �� �� �� ��   	   1      �  o BD o  g�   	   1      �  F, �4 F, ��   	   1      �  � L �  ��  �   ��   	   1      �  � �� � ��      1    , |� J �| J �| Y� |� Y� |� J      1    , (� � 8\ � 8\ �� (� �� (� �      1    , �d � � � � �� �d �� �d �      1    , �X �� � �� � � �X � �X ��   	   1      �  Q� a� Q�  u0   	   1      �   �  0�  �   ��  ܴ  ��   	   1      �  |� Q� m< Q�      1    , X �� $� �� $� �L X �L X ��   	   1      � $ �� 2� �� 2� ��  ~� ��  ~�   	   1      �  iT  �4 iT .�   	   1      �  �4  � �4 |   	   1      �  �\  g� �\ BD      1    , [� �X kH �X kH �� [� �� [� �X      1    , �( � �� � �� d �( d �( �      1    ,  d ��  ' ��  ' �  d �  d ��      1    ,  p �  ' �  ' ��  p ��  p �      1    ,  #(  �$  2�  �$  2� �  #( �  #(  �$      1    , *� �� 8\ �� 8\ � *� � *� ��      1    ,  m` 0�  }  0�  }  @P  m` @P  m` 0�   	   1      � ,  _� X  �� X  ��  ��  W�  ��  W�  �|   	   1      �  $� a� $� �L      1    , >\ �� M� �� M� �4 >\ �4 >\ ��   	   1      �  el a� el �(   	   1      �  #  �4 # .�   	   1      �   }  6�  �� 6�      1    , �� �X �t �X �t �� �� �� �� �X   	   1      �   �l s  �l ��      *    ,      � Ҩ  � Ҩ ��     ��      �             iT  � GND              iT �8 VDD               �  � R               Bh  � D              �\  � Q              q   � QB             >\  � CLK      �     � 	   0 - 
nor02     +    ,  ix  e�  S�  e�  S�  y  ix  y  ix  e� +  ,2       0    ,  c�  kl  [�  kl  [�  s<  c�  s<  c�  kl      1    ,  g�  g�  W�  g�  W�  w$  g�  w$  g�  g� +  ,1       .    ,  S�  [�  L,  [�  L,  e�  S�  e�  S�  [� +  ,3       .    ,  S�  y  L,  y  L,  ��  S�  ��  S�  y +  ,4       .    ,  S�  e�  L,  e�  L,  y  S�  y  S�  e�      0    ,  D\  kl  <�  kl  <�  s<  D\  s<  D\  kl      1    ,  HD  g�  8�  g�  8�  w$  HD  w$  HD  g� +  ,5       .    ,  4�  [�  ,�  [�  ,�  e�  4�  e�  4�  [� +  ,6       .    ,  4�  y  ,�  y  ,�  ��  4�  ��  4�  y +  ,7       .    ,  4�  e�  ,�  e�  ,�  y  4�  y  4�  e�      0    ,  %  kl  L  kl  L  s<  %  s<  %  kl      1    ,  )  g�  d  g�  d  w$  )  w$  )  g� +  ,8       +    ,  ix  e�  p  e�  p  y  ix  y  ix  e�      )    ,  ��  N       N       ��  ��  ��  ��  N  +  ,10      -    ,  qH  ]�  �  ]�  �  ��  qH  ��  qH  ]�      +    ,  ,�  e�  p  e�  p  y  ,�  y  ,�  e� +  ,9       +    ,  a� (�  L, (�  L, kH  a� kH  a� (� +  ,2       0    ,  [� .�  S� .�  S� 6�  [� 6�  [� .�      0    ,  [� F,  S� F,  S� M�  [� M�  [� F,      0    ,  [� ]�  S� ]�  S� el  [� el  [� ]�      1    ,  _� *�  P *�  P iT  _� iT  _� *� +  ,1       .    ,  L,   D\   D\ (�  L, (�  L,  +  ,3       .    ,  L, kH  D\ kH  D\ u  L, u  L, kH +  ,4       .    ,  L, (�  D\ (�  D\ kH  L, kH  L, (�      .    ,  4�   ,�   ,� (�  4� (�  4�  +  ,5       .    ,  4� kH  ,� kH  ,� u  4� u  4� kH +  ,6       .    ,  4� (�  ,� (�  ,� kH  4� kH  4� (�      0    ,  % .�  L .�  L 6�  % 6�  % .�      0    ,  % F,  L F,  L M�  % M�  % F,      0    ,  % ]�  L ]�  L el  % el  % ]�      1    ,  ) *�  d *�  d iT  ) iT  ) *� +  ,7       +    ,  a� (�  p (�  p kH  a� kH  a� (�      *    ,  y p     p     ��  y ��  y p +  ,9       ,    ,  ix !  � !  � s  ix s  ix !      +    ,  ,� (�  p (�  p kH  ,� kH  ,� (� +  ,8    
  via  �    @t  ��   
  via  �    c�  ��   
  via  �    L  ��      3    ,  6�  ��  J8  ��  J8  �`  6�  �`  6�  ��      3    ,  Y�  ��  m`  ��  m`  �`  Y�  �`  Y�  ��      3    ,  �  ��  '  ��  '  �`  �  �`  �  ��      1    ,     ��  �� ��  �� ��     ��     ��      1    ,          ��      ��  '      '              �    ,          ��      �� ��     ��              .    ,  Y�  ��  m`  ��  m`  �`  Y�  �`  Y�  ��      .    ,  �  ��  '  ��  '  �`  �  �`  �  ��   	   .      � $  0�   0�  �   #(  �   #(  �`   	   .      �   #(  ��  #(  ��  4�  ��   	   .      �   L,  ��  ]�  ��  ]�  ��   	   .      �   D\ 4  ]� 4  ]�  �`      /    ,  _�  ܴ  g�  ܴ  g�  �  _�  �  _�  ܴ      /    ,  d  ܴ  !4  ܴ  !4  �  d  �  d  ܴ      )    ,          ��      ��  ��      ��              *    ,     p  �� p  �� ��     ��     p      ,    ,  �  �  u0  �  u0  *�  �  *�  �  �      ,    ,  �  *�  2�  *�  2�  ]�  �  ]�  �  *�      ,    ,  N   *�  qH  *�  qH  ]�  N   ]�  N   *�      -    ,  � ��  u0 ��  u0 ��  � ��  � ��      -    ,  FP s  ix s  ix ��  FP ��  FP s      0    ,  0�  |  8�  |  8�  L  0�  L  0�  |      0    ,  HD  |  P  |  P  L  HD  L  HD  |      0    ,  _�  |  g�  |  g�  L  _�  L  _�  |      0    ,  d  |  !4  |  !4  L  d  L  d  |      0    ,  d �t  !4 �t  !4 �D  d �D  d �t      0    ,  0� �t  8� �t  8� �D  0� �D  0� �t      0    ,  HD �t  P �t  P �D  HD �D  HD �t      0    ,  _� �t  g� �t  g� �D  _� �D  _� �t      0    ,  [�  HD  c�  HD  c�  P  [�  P  [�  HD      0    ,  L  HD  %  HD  %  P  L  P  L  HD      0    ,  [�  0�  c�  0�  c�  8�  [�  8�  [�  0�      0    ,  L  0�  %  0�  %  8�  L  8�  L  0�      0    ,  S� �4  [� �4  [� �  S� �  S� �4      0    ,  S� ��  [� ��  [� ��  S� ��  S� ��      1    ,  [�  ��  kl  ��  kl  �l  [�  �l  [�  ��   	   1      � $  !4 *�  !4 �  @t �  @t  �`      1    ,  |  ��  %  ��  %  �l  |  �l  |  ��   	   1      �   @t  ��  @t  w$      1    ,  d  '  )  '  )  S�  d  S�  d  '      1    ,  Y�  S�  g�  S�  g�  g�  Y�  g�  Y�  S�      1    ,  d  S�  '  S�  '  g�  d  g�  d  S�      1    ,  W�  '  g�  '  g�  S�  W�  S�  W�  '      1    ,  R iT  _� iT  _� |�  R |�  R iT      1    ,  P |�  _� |�  _� ��  P ��  P |�      +    ,  �  �  m`  �  m`  #(  �  #(  �  �      +    ,  � ��  m` ��  m` �   � �   � ��      +    ,  p  U�  )  U�  )  e�  p  e�  p  U�      +    ,  p  #(  *�  #(  *�  U�  p  U�  p  #(      +    ,  W�  U�  ix  U�  ix  e�  W�  e�  W�  U�      +    ,  U�  #(  ix  #(  ix  U�  U�  U�  U�  #(      +    ,  P kH  a� kH  a� z�  P z�  P kH      +    ,  N  z�  a� z�  a� ��  N  ��  N  z�              @t  � GND  +  ,1               @t �8 VDD  +  ,1               L  �� A1 +  ,1               c�  �� A0 +  ,1               @t  �� Y  +  ,1               @t  � GND               @t �8 VDD               L  �� A1              c�  �� A0              @t  �� Y      �    , 3� 	   0 
 
inv01     +    ,  p  e�  ,�  e�  ,�  y  p  y  p  e� +  ,2       0    ,  L  kl  %  kl  %  s<  L  s<  L  kl      1    ,  d  g�  )  g�  )  w$  d  w$  d  g� +  ,1       .    ,  ,�  [�  4�  [�  4�  e�  ,�  e�  ,�  [� +  ,3       .    ,  ,�  y  4�  y  4�  ��  ,�  ��  ,�  y +  ,4       .    ,  ,�  e�  4�  e�  4�  y  ,�  y  ,�  e�      0    ,  <�  kl  D\  kl  D\  s<  <�  s<  <�  kl      1    ,  8�  g�  HD  g�  HD  w$  8�  w$  8�  g� +  ,5       +    ,  p  e�  J8  e�  J8  y  p  y  p  e�      )    ,      N   a�  N   a�  ��      ��      N  +  ,7       -    ,  �  ]�  R  ]�  R  ��  �  ��  �  ]�      +    ,  4�  e�  J8  e�  J8  y  4�  y  4�  e� +  ,6       +    ,  p 8�  ,� 8�  ,� cx  p cx  p 8� +  ,2       0    ,  L >\  % >\  % F,  L F,  L >\      0    ,  L U�  % U�  % ]�  L ]�  L U�      1    ,  d :t  ) :t  ) a�  d a�  d :t +  ,1       .    ,  ,� .�  4� .�  4� 8�  ,� 8�  ,� .� +  ,3       .    ,  ,� cx  4� cx  4� m<  ,� m<  ,� cx +  ,4       .    ,  ,� 8�  4� 8�  4� cx  ,� cx  ,� 8�      0    ,  <� >\  D\ >\  D\ F,  <� F,  <� >\      0    ,  <� U�  D\ U�  D\ ]�  <� ]�  <� U�      1    ,  8� :t  HD :t  HD a�  8� a�  8� :t +  ,5       +    ,  p 8�  J8 8�  J8 cx  p cx  p 8�      *    ,     !  a� !  a� z�     z�     ! +  ,7       ,    ,  � 0�  R 0�  R kH  � kH  � 0�      +    ,  4� 8�  J8 8�  J8 cx  4� cx  4� 8� +  ,6    
  via    '  �   
  via    J8  �      1    ,          a�      a�  '      '              1    ,     ��  a� ��  a� ��     ��     ��      1    ,          a�      a�  '      '              1    ,     ��  a� ��  a� ��     ��     ��      3    ,  L  �P  0�  �P  0�  ��  L  ��  L  �P      3    ,  @t  �P  S�  �P  S�  ��  @t  ��  @t  �P      �    ,          a�      a� ��     ��              �    ,  !4  �D  0�  �D  0�  ��  !4  ��  !4  �D      /    ,  %  �,  ,�  �,  ,�  ��  %  ��  %  �,   	   .      �   0� .�  0�  ��      .    ,  @  �P  2�  �P  2�  ��  @  ��  @  �P      )    ,          a�      a�  ��      ��              *    ,     !  a� !  a� ��     ��     !      -    ,  � ��  Y� ��  Y� ��  � ��  � ��      -    ,  � kH  2� kH  2� ��  � ��  � kH      ,    ,  �  �  Y�  �  Y�  *�  �  *�  �  �      ,    ,  �  *�  2�  *�  2�  ]�  �  ]�  �  *�      +    ,  �  �  R  �  R  #(  �  #(  �  �      +    ,  � ��  R ��  R �   � �   � ��      +    ,  p s  *� s  *� ��  p ��  p s      +    ,  p cx  ) cx  ) s  p s  p cx      +    ,  p  U�  )  U�  )  e�  p  e�  p  U�      +    ,  p  #(  *�  #(  *�  U�  p  U�  p  #(   	   1      �   Bh :t  Bh  w$      1    ,  !4  �D  0�  �D  0�  ��  !4  ��  !4  �D      1    ,  d a�  ' a�  ' u  d u  d a�      1    ,  d u  ) u  ) ��  d ��  d u      1    ,  d  S�  '  S�  '  g�  d  g�  d  S�      1    ,  d  '  )  '  )  S�  d  S�  d  '      0    ,  D\  |  L,  |  L,  L  D\  L  D\  |      0    ,  ,�  |  4�  |  4�  L  ,�  L  ,�  |      0    ,  |  |  L  |  L  L  |  L  |  |      0    ,  D\ �t  L, �t  L, �D  D\ �D  D\ �t      0    ,  ,� �t  4� �t  4� �D  ,� �D  ,� �t      0    ,  | �t  L �t  L �D  | �D  | �t      0    ,  L x�  % x�  % ��  L ��  L x�      0    ,  L �d  % �d  % �4  L �4  L �d      0    ,  L  HD  %  HD  %  P  L  P  L  HD      0    ,  L  0�  %  0�  %  8�  L  8�  L  0�              0�  � GND  +  ,1               0� �8 VDD  +  ,1               J8  � Y  +  ,1               '  � A  +  ,1               0�  � GND               0� �8 VDD               J8  � Y               '  � A      �   
  ,� 	   /  
aoi32     0    ,  L BD  % BD  % J  L J  L BD      0    ,  L Y�  % Y�  % a�  L a�  L Y�      0    ,  L q$  % q$  % x�  L x�  L q$      1    ,  d >\  ) >\  ) |�  d |�  d >\ +  ,1       .    ,  ,� 2�  4� 2�  4� <h  ,� <h  ,� 2� +  ,3       .    ,  ,� ~�  4� ~�  4� ��  ,� ��  ,� ~� +  ,4       .    ,  ,� <h  4� <h  4� ~�  ,� ~�  ,� <h      0    ,  <� BD  D\ BD  D\ J  <� J  <� BD      0    ,  <� Y�  D\ Y�  D\ a�  <� a�  <� Y�      0    ,  <� q$  D\ q$  D\ x�  <� x�  <� q$      1    ,  8� >\  HD >\  HD |�  8� |�  8� >\ +  ,5       .    ,  L, 2�  S� 2�  S� <h  L, <h  L, 2� +  ,6       .    ,  L, ~�  S� ~�  S� ��  L, ��  L, ~� +  ,7       .    ,  L, <h  S� <h  S� ~�  L, ~�  L, <h      0    ,  [� BD  c� BD  c� J  [� J  [� BD      0    ,  [� Y�  c� Y�  c� a�  [� a�  [� Y�      0    ,  [� q$  c� q$  c� x�  [� x�  [� q$      1    ,  W� >\  g� >\  g� |�  W� |�  W� >\ +  ,8       .    ,  kl 2�  s< 2�  s< <h  kl <h  kl 2� +  ,9       .    ,  kl ~�  s< ~�  s< ��  kl ��  kl ~� +  ,10      .    ,  kl <h  s< <h  s< ~�  kl ~�  kl <h      0    ,  { BD  �� BD  �� J  { J  { BD      0    ,  { Y�  �� Y�  �� a�  { a�  { Y�      0    ,  { q$  �� q$  �� x�  { x�  { q$      1    ,  w$ >\  �� >\  �� |�  w$ |�  w$ >\ +  ,11      .    ,  �� 2�  �| 2�  �| <h  �� <h  �� 2� +  ,12      .    ,  �� ~�  �| ~�  �| ��  �� ��  �� ~� +  ,13      .    ,  �� <h  �| <h  �| ~�  �� ~�  �� <h      0    ,  �L BD  � BD  � J  �L J  �L BD      0    ,  �L Y�  � Y�  � a�  �L a�  �L Y�      0    ,  �L q$  � q$  � x�  �L x�  �L q$      1    ,  �d >\  � >\  � |�  �d |�  �d >\ +  ,14      .    ,  �� 2�  �� 2�  �� <h  �� <h  �� 2� +  ,15      .    ,  �� ~�  �� ~�  �� ��  �� ��  �� ~� +  ,16      .    ,  �� <h  �� <h  �� ~�  �� ~�  �� <h      0    ,  �� BD  �\ BD  �\ J  �� J  �� BD      0    ,  �� Y�  �\ Y�  �\ a�  �� a�  �� Y�      0    ,  �� q$  �\ q$  �\ x�  �� x�  �� q$      1    ,  �� >\  �D >\  �D |�  �� |�  �� >\ +  ,17      +    ,  p <h  �8 <h  �8 ~�  p ~�  p <h      *    ,     $�  ި $�  ި �@     �@     $� +  ,19      ,    ,  � 4�  � 4�  � ��  � ��  � 4�      +    ,  p <h  ,� <h  ,� ~�  p ~�  p <h +  ,2       +    ,  �� <h  �8 <h  �8 ~�  �� ~�  �� <h +  ,18      +    ,  p  L,  ,�  L,  ,�  ��  p  ��  p  L, +  ,2       0    ,  L  R  %  R  %  Y�  L  Y�  L  R      0    ,  L  ix  %  ix  %  qH  L  qH  L  ix      0    ,  L  ��  %  ��  %  ��  L  ��  L  ��      1    ,  d  N   )  N   )  ��  d  ��  d  N  +  ,1       .    ,  ,�  Bh  4�  Bh  4�  L,  ,�  L,  ,�  Bh +  ,3       .    ,  ,�  ��  4�  ��  4�  �X  ,�  �X  ,�  �� +  ,4       .    ,  ,�  L,  4�  L,  4�  ��  ,�  ��  ,�  L,      .    ,  D\  Bh  L,  Bh  L,  L,  D\  L,  D\  Bh +  ,5       .    ,  D\  ��  L,  ��  L,  �X  D\  �X  D\  �� +  ,6       .    ,  D\  L,  L,  L,  L,  ��  D\  ��  D\  L,      .    ,  [�  Bh  c�  Bh  c�  L,  [�  L,  [�  Bh +  ,7       .    ,  [�  ��  c�  ��  c�  �X  [�  �X  [�  �� +  ,8       .    ,  [�  L,  c�  L,  c�  ��  [�  ��  [�  L,      0    ,  kl  R  s<  R  s<  Y�  kl  Y�  kl  R      0    ,  kl  ix  s<  ix  s<  qH  kl  qH  kl  ix      0    ,  kl  ��  s<  ��  s<  ��  kl  ��  kl  ��      1    ,  g�  N   w$  N   w$  ��  g�  ��  g�  N  +  ,9       .    ,  }   Y�  ��  Y�  ��  c�  }   c�  }   Y� +  ,10      .    ,  }   ��  ��  ��  ��  �X  }   �X  }   �� +  ,11      .    ,  }   c�  ��  c�  ��  ��  }   ��  }   c�      .    ,  �p  Y�  �@  Y�  �@  c�  �p  c�  �p  Y� +  ,12      .    ,  �p  ��  �@  ��  �@  �X  �p  �X  �p  �� +  ,13      .    ,  �p  c�  �@  c�  �@  ��  �p  ��  �p  c�      0    ,  �  ix  ��  ix  ��  qH  �  qH  �  ix      0    ,  �  ��  ��  ��  ��  ��  �  ��  �  ��      1    ,  �(  e�  ��  e�  ��  ��  �(  ��  �(  e� +  ,14      +    <  y  L,  y  c�  ��  c�  ��  ��  p  ��  p  L,  y  L,      )    <  ��  4�  ��  L,  �,  L,  �,  �      �      4�  ��  4� +  ,16      -    <  ��  D\  ��  [�  ��  [�  ��  �d  �  �d  �  D\  ��  D\      +    ,  �@  c�  ��  c�  ��  ��  �@  ��  �@  c� +  ,15   
  via  �  B�         8�  �   
  via  �  B�         ~�  �   
  via  �  B�         �D  �   
  via  �  B�         �  �   
  via  �  B�         [�  �   
  via  �  B�         |  �      3    ,  �X  �P  ��  �P  ��  ��  �X  ��  �X  �P      3    ,  ��  �P  �  �P  �  ��  ��  ��  ��  �P      3    ,  �  �P  @  �P  @  ��  �  ��  �  �P      3    ,  .�  �P  Bh  �P  Bh  ��  .�  ��  .�  �P      3    ,  R  �P  e�  �P  e�  ��  R  ��  R  �P      3    ,  u0  �P  ��  �P  ��  ��  u0  ��  u0  �P      1    ,     ��  ި ��  ި ��     ��     ��      1    ,          ި      ި  '      '              0    ,  0�  |  8�  |  8�  L  0�  L  0�  |      0    ,  HD  |  P  |  P  L  HD  L  HD  |      0    ,  _�  |  g�  |  g�  L  _�  L  _�  |      0    ,  w$  |  ~�  |  ~�  L  w$  L  w$  |      0    ,  ��  |  �d  |  �d  L  ��  L  ��  |      0    ,  �  |  ��  |  ��  L  �  L  �  |      0    ,  �t  |  �D  |  �D  L  �t  L  �t  |      0    ,  d  |  !4  |  !4  L  d  L  d  |      0    ,  w$ �t  ~� �t  ~� �D  w$ �D  w$ �t      0    ,  _� �t  g� �t  g� �D  _� �D  _� �t      0    ,  HD �t  P �t  P �D  HD �D  HD �t      0    ,  0� �t  8� �t  8� �D  0� �D  0� �t      0    ,  �� �t  �d �t  �d �D  �� �D  �� �t      0    ,  � �t  �� �t  �� �D  � �D  � �t      0    ,  �t �t  �D �t  �D �D  �t �D  �t �t      0    ,  d �t  !4 �t  !4 �D  d �D  d �t      0    ,  L �L  % �L  % �  L �  L �L      0    ,  [� �L  c� �L  c� �  [� �  [� �L      0    ,  L  .�  %  .�  %  6�  L  6�  L  .�      0    ,  �  FP  ��  FP  ��  N   �  N   �  FP      0    ,  �  .�  ��  .�  ��  6�  �  6�  �  .�   	   1      � $  �� |�  �� �@  �� �@  �� |�   	   1      � $  �@ >\  �@ d  ~� d  ~�  ��      1    ,  �  R  ��  R  ��  e�  �  e�  �  R   	   1      � $  qH  ��  qH  ��  {  ��  {  �P   	   1      � $  }  >\  }  *�  Bh *�  Bh >\      1    ,  �(  '  ��  '  ��  R  �(  R  �(  '      1    ,  S�  �D  c�  �D  c�  ��  S�  ��  S�  �D      1    ,  �L  �D  ��  �D  ��  ��  �L  ��  �L  �D      1    ,  �  �D  L  �D  L  ��  �  ��  �  �D      1    ,  0�  �D  @t  �D  @t  ��  0�  ��  0�  �D      1    ,  �t  �D  �  �D  �  ��  �t  ��  �t  �D      1    ,  d |�  ' |�  ' �d  d �d  d |�      1    ,  d �d  ) �d  ) ��  d ��  d �d      1    ,  W� �d  g� �d  g� ��  W� ��  W� �d      1    ,  Y� |�  e� |�  e� �d  Y� �d  Y� |�      1    ,  d  :�  '  :�  '  N   d  N   d  :�      1    ,  d  '  )  '  )  :�  d  :�  d  '      +    ,  �  �  �   �  �   #(  �  #(  �  �      +    ,  � ��  �  ��  �  �   � �   � ��      +    ,  p ~�  ) ~�  ) �p  p �p  p ~�      +    ,  p �p  *� �p  *� ��  p ��  p �p      +    ,  U� �p  ix �p  ix ��  U� ��  U� �p      +    ,  W� ~�  g� ~�  g� �p  W� �p  W� ~�      +    ,  p  <�  )  <�  )  L,  p  L,  p  <�      +    ,  p  #(  *�  #(  *�  <�  p  <�  p  #(      +    ,  �(  S�  ��  S�  ��  c�  �(  c�  �(  S�      +    ,  �4  #(  ��  #(  ��  S�  �4  S�  �4  #(      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      ,    ,  �  *�  2�  *�  2�  D\  �  D\  �  *�      ,    ,  �d  *�  ��  *�  ��  [�  �d  [�  �d  *�      -    ,  � ��  �� ��  �� ��  � ��  � ��      -    ,  � ��  2� ��  2� ��  � ��  � ��      -    ,  N  ��  qH ��  qH ��  N  ��  N  ��      )    ,          ި      ި  �      �              *    ,     $�  ި $�  ި ��     ��     $�      /    ,  W�  �,  _�  �,  _�  ��  W�  ��  W�  �,      /    ,  �4  �,  �  �,  �  ��  �4  ��  �4  �,      /    ,  �  �,  d  �,  d  ��  �  ��  �  �,      /    ,  4�  �,  <�  �,  <�  ��  4�  ��  4�  �,      /    ,  �\  �,  �,  �,  �,  ��  �\  ��  �\  �,   	   .      � $  >�  ��  >� (  P (  P 2�      .    ,  �  �P  @  �P  @  ��  �  ��  �  �P   	   .      � $  oT 2�  oT 	�  _� 	�  _�  �X      .    ,  �X  �P  ��  �P  ��  ��  �X  ��  �X  �P      .    ,  ��  �P  �  �P  �  ��  ��  ��  ��  �P      .    ,  R  �P  e�  �P  e�  ��  R  ��  R  �P   	   .      �   �h  �P  �h  �X  �p  �X      .    ,  .�  �P  Bh  �P  Bh  ��  .�  ��  .�  �P   	   .      �   4� 2�  X 2�  X  ��   	   .      �   X  �P  X  �X  4�  �X   	   .      � $  HD  �X  HD  ��  >�  ��  >�  �P   	   .      � $  ��  �X  ��  ��  �@  ��  �@  �P   	   .      � $  �� 2�  �� $�  �h $�  �h  ��   	   .      � $  �� 2�  �� �  �@ �  �@  ��              oT  � GND  +  ,1               oT �8 VDD  +  ,1               �  � B0 +  ,1               �D  � B1 +  ,1               |  � A2 +  ,1               8�  � A1 +  ,1               [�  � A0 +  ,1               ~�  � Y  +  ,1       �    ,          ި      ި ��     ��                      oT  � GND               oT �8 VDD               �  � B0              �D  � B1              |  � A2              8�  � A1              [�  � A0              ~�  � Y      �     	� 	   0 # 
nand02    +    <  S� O�  S� ��  ix ��  ix _�  c� _�  c� O�  S� O� +  ,2       0    ,  c� el  [� el  [� m<  c� m<  c� el      0    ,  c� |�  [� |�  [� ��  c� ��  c� |�      1    ,  g� a�  W� a�  W� ��  g� ��  g� a� +  ,1       .    ,  S� F,  L, F,  L, O�  S� O�  S� F, +  ,3       .    ,  S� ��  L, ��  L, �L  S� �L  S� �� +  ,4       .    ,  S� O�  L, O�  L, ��  S� ��  S� O�      0    ,  D\ U�  <� U�  <� ]�  D\ ]�  D\ U�      0    ,  D\ m<  <� m<  <� u  D\ u  D\ m<      1    ,  HD Q�  8� Q�  8� x�  HD x�  HD Q� +  ,5       .    ,  4� F,  ,� F,  ,� O�  4� O�  4� F, +  ,6       .    ,  4� ��  ,� ��  ,� �L  4� �L  4� �� +  ,7       .    ,  4� O�  ,� O�  ,� ��  4� ��  4� O�      0    ,  % el  L el  L m<  % m<  % el      0    ,  % |�  L |�  L ��  % ��  % |�      1    ,  ) a�  d a�  d ��  ) ��  ) a� +  ,8       +    L  L O�  L _�  p _�  p ��  ix ��  ix _�  c� _�  c� O�  L O�      *    L  � 8�  � H      H      ��  �� ��  �� H   { H   { 8�  � 8� +  ,10      ,    L  | H   | W�  � W�  � �X  qH �X  qH W�  kl W�  kl H   | H       +    <  L O�  L _�  p _�  p ��  ,� ��  ,� O�  L O� +  ,9       +    ,  p  J8  ,�  J8  ,�  u0  p  u0  p  J8 +  ,2       0    ,  L  P  %  P  %  W�  L  W�  L  P      0    ,  L  g�  %  g�  %  oT  L  oT  L  g�      1    ,  d  L,  )  L,  )  s<  d  s<  d  L, +  ,1       .    ,  ,�  @t  4�  @t  4�  J8  ,�  J8  ,�  @t +  ,3       .    ,  ,�  u0  4�  u0  4�  ~�  ,�  ~�  ,�  u0 +  ,4       .    ,  ,�  J8  4�  J8  4�  u0  ,�  u0  ,�  J8      .    ,  D\  @t  L,  @t  L,  J8  D\  J8  D\  @t +  ,5       .    ,  D\  u0  L,  u0  L,  ~�  D\  ~�  D\  u0 +  ,6       .    ,  D\  J8  L,  J8  L,  u0  D\  u0  D\  J8      0    ,  S�  P  [�  P  [�  W�  S�  W�  S�  P      0    ,  S�  g�  [�  g�  [�  oT  S�  oT  S�  g�      1    ,  P  L,  _�  L,  _�  s<  P  s<  P  L, +  ,7       +    ,  p  J8  a�  J8  a�  u0  p  u0  p  J8      )    ,      2�  y  2�  y  ��      ��      2� +  ,9       -    ,  �  Bh  ix  Bh  ix  }   �  }   �  Bh      +    ,  L,  J8  a�  J8  a�  u0  L,  u0  L,  J8 +  ,8    
  via    D\  �   
  via    !4  �   
  via    g�  �      3    ,  :�  �P  N   �P  N   ��  :�  ��  :�  �P      3    ,  ]�  �P  qH  �P  qH  ��  ]�  ��  ]�  �P      3    ,  p  �P  *�  �P  *�  ��  p  ��  p  �P      1    ,     ��  �� ��  �� ��     ��     ��      1    ,          ��      ��  '      '              1    ,     ��  �� ��  �� ��     ��     ��      1    ,          ��      ��  '      '              �    ,          ��      �� ��     ��              1    ,  <�  �D  L,  �D  L,  ��  <�  ��  <�  �D      1    ,  d  �D  )  �D  )  ��  d  ��  d  �D      1    ,  d  '  )  '  )  8�  d  8�  d  '      1    ,  d �  ) �  ) ��  d ��  d �      1    ,  d ��  ' ��  ' �  d �  d ��      1    ,  W� �  g� �  g� ��  W� ��  W� �   	   1      � $  @t Q�  @t ,�  c� ,�  c�  ��      1    ,  Y� ��  g� ��  g� �  Y� �  Y� ��      1    ,  d  8�  '  8�  '  L,  d  L,  d  8�   	   1      �   c�  �P  c�  g�      .    ,  :�  �P  N   �P  N   ��  :�  ��  :�  �P      .    ,  p  �P  *�  �P  *�  ��  p  ��  p  �P   	   .      � $  P F,  P p  J8 p  J8  ��   	   .      �   '  �P  '  ��  4�  ��   	   .      �   4� BD  ' BD  '  ��   	   .      �   HD  ~�  HD  �P      )    ,          ��      ��  ��      ��              ,    ,  �  �  u0  �  u0  *�  �  *�  �  �      ,    ,  �  *�  2�  *�  2�  Bh  �  Bh  �  *�      +    ,  �  �  m`  �  m`  #(  �  #(  �  �      +    ,  � ��  m` ��  m` �   � �   � ��      +    ,  p ��  ) ��  ) �(  p �(  p ��      +    ,  W� ��  ix ��  ix �(  W� �(  W� ��      +    ,  U� �(  ix �(  ix ��  U� ��  U� �(      +    ,  p �(  *� �(  *� ��  p ��  p �(      +    ,  p  :�  )  :�  )  J8  p  J8  p  :�      +    ,  p  #(  *�  #(  *�  :�  p  :�  p  #(      0    ,  0�  |  8�  |  8�  L  0�  L  0�  |      0    ,  HD  |  P  |  P  L  HD  L  HD  |      0    ,  _�  |  g�  |  g�  L  _�  L  _�  |      0    ,  d  |  !4  |  !4  L  d  L  d  |      0    ,  d �t  !4 �t  !4 �D  d �D  d �t      0    ,  0� �t  8� �t  8� �D  0� �D  0� �t      0    ,  HD �t  P �t  P �D  HD �D  HD �t      0    ,  _� �t  g� �t  g� �D  _� �D  _� �t      0    ,  [� �  c� �  c� ��  [� ��  [� �      0    ,  L �  % �  % ��  L ��  L �      0    ,  L  ,�  %  ,�  %  4�  L  4�  L  ,�      *    ,     8�  �� 8�  �� ��     ��     8�      -    ,  � ��  u0 ��  u0 ��  � ��  � ��      -    ,  � �X  2� �X  2� ��  � ��  � �X      -    ,  N  �X  qH �X  qH ��  N  ��  N  �X      /    ,  @t  �,  HD  �,  HD  ��  @t  ��  @t  �,      /    ,  L  �,  %  �,  %  ��  L  ��  L  �,              @t  � GND  +  ,1               @t �8 VDD  +  ,1               !4  � A1 +  ,1               D\  � A0 +  ,1               g�  � Y  +  ,1               @t  � GND               @t �8 VDD               !4  � A1              D\  � A0              g�  � Y      �     +� 	   0  
mux21     +    ,  p  ]�  ,�  ]�  ,�  ��  p  ��  p  ]� +  ,2       0    ,  L  c�  %  c�  %  kl  L  kl  L  c�      0    ,  L  {  %  {  %  ��  L  ��  L  {      1    ,  d  _�  )  _�  )  ��  d  ��  d  _� +  ,1       .    ,  ,�  S�  4�  S�  4�  ]�  ,�  ]�  ,�  S� +  ,3       .    ,  ,�  ��  4�  ��  4�  �|  ,�  �|  ,�  �� +  ,4       .    ,  ,�  ]�  4�  ]�  4�  ��  ,�  ��  ,�  ]�      .    ,  D\  S�  L,  S�  L,  ]�  D\  ]�  D\  S� +  ,5       .    ,  D\  ��  L,  ��  L,  �|  D\  �|  D\  �� +  ,6       .    ,  D\  ]�  L,  ]�  L,  ��  D\  ��  D\  ]�      0    ,  S�  c�  [�  c�  [�  kl  S�  kl  S�  c�      0    ,  S�  {  [�  {  [�  ��  S�  ��  S�  {      1    ,  P  _�  _�  _�  _�  ��  P  ��  P  _� +  ,7       .    ,  c�  S�  kl  S�  kl  ]�  c�  ]�  c�  S� +  ,8       .    ,  c�  ��  kl  ��  kl  �|  c�  �|  c�  �� +  ,9       .    ,  c�  ]�  kl  ]�  kl  ��  c�  ��  c�  ]�      .    ,  {  S�  ��  S�  ��  ]�  {  ]�  {  S� +  ,10      .    ,  {  ��  ��  ��  ��  �|  {  �|  {  �� +  ,11      .    ,  {  ]�  ��  ]�  ��  ��  {  ��  {  ]�      0    ,  ��  c�  �|  c�  �|  kl  ��  kl  ��  c�      0    ,  ��  {  �|  {  �|  ��  ��  ��  ��  {      1    ,  ��  _�  �d  _�  �d  ��  ��  ��  ��  _� +  ,12      .    ,  �@  kl  �  kl  �  u0  �@  u0  �@  kl +  ,13      .    ,  �@  ��  �  ��  �  �|  �@  �|  �@  �� +  ,14      .    ,  �@  u0  �  u0  �  ��  �@  ��  �@  u0      0    ,  ��  {  ��  {  ��  ��  ��  ��  ��  {      1    ,  ��  w$  ��  w$  ��  ��  ��  ��  ��  w$ +  ,15      +    <  �X  ]�  �X  u0  ��  u0  ��  ��  p  ��  p  ]�  �X  ]�      )    <  ��  FP  ��  ]�  ��  ]�  ��  �(      �(      FP  ��  FP +  ,17      -    <  �(  U�  �(  m`  �\  m`  �\  ��  �  ��  �  U�  �(  U�      +    ,  �  u0  ��  u0  ��  ��  �  ��  �  u0 +  ,16      0    ,  L 6�  % 6�  % >\  L >\  L 6�      0    ,  L M�  % M�  % U�  L U�  L M�      0    ,  L el  % el  % m<  L m<  L el      1    ,  d 2�  ) 2�  ) q$  d q$  d 2� +  ,1       .    ,  ,� d  4� d  4� (  ,� (  ,� d +  ,3       .    ,  ,� s  4� s  4� |�  ,� |�  ,� s +  ,4       .    ,  ,� (  4� (  4� s  ,� s  ,� (      .    ,  D\ d  L, d  L, (  D\ (  D\ d +  ,5       .    ,  D\ s  L, s  L, |�  D\ |�  D\ s +  ,6       .    ,  D\ (  L, (  L, s  D\ s  D\ (      0    ,  S� #  [� #  [� *�  S� *�  S� #      0    ,  S� :t  [� :t  [� BD  S� BD  S� :t      0    ,  S� Q�  [� Q�  [� Y�  S� Y�  S� Q�      1    ,  P   _�   _� ]�  P ]�  P  +  ,7       .    ,  c� d  kl d  kl (  c� (  c� d +  ,8       .    ,  c� s  kl s  kl |�  c� |�  c� s +  ,9       .    ,  c� (  kl (  kl s  c� s  c� (      .    ,  { d  �� d  �� (  { (  { d +  ,10      .    ,  { s  �� s  �� |�  { |�  { s +  ,11      .    ,  { (  �� (  �� s  { s  { (      0    ,  �� 6�  �| 6�  �| >\  �� >\  �� 6�      0    ,  �� M�  �| M�  �| U�  �� U�  �� M�      0    ,  �� el  �| el  �| m<  �� m<  �� el      1    ,  �� 2�  �d 2�  �d q$  �� q$  �� 2� +  ,12      .    ,  �@ d  � d  � (  �@ (  �@ d +  ,13      .    ,  �@ H   � H   � Q�  �@ Q�  �@ H  +  ,14      .    ,  �@ (  � (  � H   �@ H   �@ (      0    ,  �� #  �� #  �� *�  �� *�  �� #      0    ,  �� :t  �� :t  �� BD  �� BD  �� :t      1    ,  ��   ��   �� F,  �� F,  ��  +  ,15      +    L  �� (  �� H   �X H   �X s  p s  p 0�  L 0�  L (  �� (      *    L  �� �  �� _�  �� _�  �� ��     ��     @  � @  � �  �� � +  ,17      ,    L  �\ X  �\ O�  �( O�  �( z�  � z�  � (�  | (�  | X  �\ X      +    <  ,� (  ,� s  p s  p 0�  L 0�  L (  ,� ( +  ,2       +    ,  � (  �� (  �� H   � H   � ( +  ,16   
  via  �  B�         �L  �   
  via    m`  �   
  via    L  �   
  via    J8  �      3    ,  ��  �P  �  �P  �  ��  ��  ��  ��  �P      3    ,  �  �P  '  �P  '  ��  �  ��  �  �P      3    ,  c�  �P  w$  �P  w$  ��  c�  ��  c�  �P      3    ,  @t  �P  S�  �P  S�  ��  @t  ��  @t  �P      1    ,          ��      ��  '      '              1    ,     ��  �� ��  �� ��     ��     ��      �    ,          ��      �� ��     ��              1    ,  e�  �D  u0  �D  u0  ��  e�  ��  e�  �D      1    ,  d q$  ' q$  ' ��  d ��  d q$      1    ,  �|  �D  �  �D  �  ��  �|  ��  �|  �D      1    ,  {  �H  ��  �H  ��  ��  {  ��  {  �H   	   1      � $  !4  �P  !4  �(  W�  �(  W�  ��      1    ,  d ��  ) ��  ) ��  d ��  d ��      1    ,  p  '  '  '  '  L,  p  L,  p  '      1    ,  ��  '  �p  '  �p  >�  ��  >�  ��  '      1    ,  Bh  �D  R  �D  R  ��  Bh  ��  Bh  �D      1    ,  ��  >�  �d  >�  �d  N   ��  N   ��  >�   	   1      �   ��  {  �� *�   	   1      �   {  �$  N   �$  N   ��   	   1      � $  U�   U� �  !4 �  !4  ��      1    ,  d  L,  '  L,  '  _�  d  _�  d  L,   	   1      �   ��  w$  ��  Bh      1    ,  ��  N   �d  N   �d  _�  ��  _�  ��  N       1    ,  �  2�  ��  2�  ��  Bh  �  Bh  �  2�      1    ,  �� ��  �d ��  �d ��  �� ��  �� ��      1    ,  �� q$  �d q$  �d ��  �� ��  �� q$      +    ,  p ��  �� ��  �� �   p �   p ��      +    ,  |  �  ��  �  ��  #(  |  #(  |  �      +    ,  |  #(  )  #(  )  N   |  N   |  #(      +    ,  p  N   )  N   )  ]�  p  ]�  p  N       +    ,  ��  <�  �X  <�  �X  P  ��  P  ��  <�      +    ,  p ��  *� ��  *� ��  p ��  p ��      +    ,  �� ��  �X ��  �X ��  �� ��  �� ��      +    ,  �� s  �X s  �X ��  �� ��  �� s      +    ,  p s  ) s  ) ��  p ��  p s      +    ,  ��  P  �X  P  �X  ]�  ��  ]�  ��  P      0    ,  L  |  %  |  %  L  L  L  L  |      0    ,  4�  |  <�  |  <�  L  4�  L  4�  |      0    ,  c�  |  kl  |  kl  L  c�  L  c�  |      0    ,  L,  |  S�  |  S�  L  L,  L  L,  |      0    ,  {  |  ��  |  ��  L  {  L  {  |      0    ,  �| �t  �L �t  �L �D  �| �D  �| �t      0    ,  �|  |  �L  |  �L  L  �|  L  �|  |      0    ,  { �t  �� �t  �� �D  { �D  { �t      0    ,  ��  |  ��  |  ��  L  ��  L  ��  |      0    ,  L �t  % �t  % �D  L �D  L �t      0    ,  4� �t  <� �t  <� �D  4� �D  4� �t      0    ,  L, �t  S� �t  S� �D  L, �D  L, �t      0    ,  c� �t  kl �t  kl �D  c� �D  c� �t      0    ,  �� �t  �� �t  �� �D  �� �D  �� �t      0    ,  X  >�  #(  >�  #(  FP  X  FP  X  >�      0    ,  L ��  % ��  % �d  L �d  L ��      0    ,  �� ��  �| ��  �| �d  �� �d  �� ��      0    ,  �� �  �| �  �| ��  �� ��  �� �      0    ,  L �  % �  % ��  L ��  L �      0    ,  ��  Bh  �|  Bh  �|  J8  ��  J8  ��  Bh      .    ,  c�  �P  w$  �P  w$  ��  c�  ��  c�  �P   	   .      �   HD  �|  HD  �P      .    ,  ��  �P  �  �P  �  ��  ��  ��  ��  �P   	   .      �   0� d  0�  �|   	   .      �   {  �d  �@  �d   	   .      �   g� d  g�  ��  y  ��   	   .      � $  g�  ��  g�  �x  HD  �x  HD d   	   .      �   g�  �|  g�  �P      .    ,  @t  �P  S�  �P  S�  ��  @t  ��  @t  �P   	   .      �   { |  �@ |   	   .      �   �( d  �(  �|      .    ,  y  �T  ��  �T  ��  ��  y  ��  y  �T      .    ,  �  0�  ��  0�  ��  D\  �  D\  �  0�   	   .      �   0�  S�  0�  4�  �  4�      /    ,  �d  �,  �4  �,  �4  ��  �d  ��  �d  �,      /    ,  ix  �,  qH  �,  qH  ��  ix  ��  ix  �,      /    ,  FP  �,  N   �,  N   ��  FP  ��  FP  �,      /    ,  ~�  �0  ��  �0  ��  �   ~�  �   ~�  �0      /    ,  ��  6�  ��  6�  ��  >�  ��  >�  ��  6�      -    ,  � ��  �h ��  �h ��  � ��  � ��      -    ,  � z�  2� z�  2� ��  � ��  � z�      -    ,  }  z�  �( z�  �( ��  }  ��  }  z�      )    ,          ��      ��  �(      �(              *    ,     �  �� �  �� ��     ��     �      ,    ,  �  *�  0�  *�  0�  U�  �  U�  �  *�      ,    ,  �  �  �h  �  �h  *�  �  *�  �  �      ,    ,  }   *�  �(  *�  �(  U�  }   U�  }   *�              h~  � GND  +  ,1               h~ �8 VDD  +  ,1               L  � Y  +  ,1               �L  � S0 +  ,1               m`  � A1 +  ,1               J8  � A0 +  ,1               h~  � GND               h~ �8 VDD               L  � Y               �L  � S0              m`  � A1              J8  � A0     �   	 4 � 	   "  nor02ii     +    ,  p @  ,� @  ,� D8  p D8  p @ +  ,2       0    ,  L   %   % &�  L &�  L       0    ,  L 6�  % 6�  % >\  L >\  L 6�      1    ,  d 4  ) 4  ) BD  d BD  d 4 +  ,1       .    ,  ,� |  4� |  4� @  ,� @  ,� | +  ,3       .    ,  ,� D8  4� D8  4� M�  ,� M�  ,� D8 +  ,4       .    ,  ,� @  4� @  4� D8  ,� D8  ,� @      0    ,  >�   FP   FP &�  >� &�  >�       0    ,  >� 6�  FP 6�  FP >\  >� >\  >� 6�      0    ,  >� M�  FP M�  FP U�  >� U�  >� M�      1    ,  :� 4  J8 4  J8 Y�  :� Y�  :� 4 +  ,5       .    ,  N  |  U� |  U� @  N  @  N  | +  ,6       .    ,  N  [�  U� [�  U� el  N  el  N  [� +  ,7       .    ,  N  @  U� @  U� [�  N  [�  N  @      .    ,  e� |  m` |  m` @  e� @  e� | +  ,8       .    ,  e� [�  m` [�  m` el  e� el  e� [� +  ,9       .    ,  e� @  m` @  m` [�  e� [�  e� @      0    ,  u0   }    }  &�  u0 &�  u0       0    ,  u0 6�  }  6�  }  >\  u0 >\  u0 6�      0    ,  u0 M�  }  M�  }  U�  u0 U�  u0 M�      1    ,  qH 4  �� 4  �� Y�  qH Y�  qH 4 +  ,10      +    <  �� @  �� [�  8� [�  8� D8  p D8  p @  �� @      *    <  �L �  �L s  !4 s  !4 [�     [�     �  �L � +  ,12      ,    <  �� p  �� cx  0� cx  0� L  � L  � p  �� p      +    ,  m` @  �� @  �� [�  m` [�  m` @ +  ,11      +    ,  ��  e�  s<  e�  s<  y  ��  y  ��  e� +  ,2       0    ,  ��  kl  {  kl  {  s<  ��  s<  ��  kl      1    ,  ��  g�  w$  g�  w$  w$  ��  w$  ��  g� +  ,1       .    ,  s<  [�  kl  [�  kl  e�  s<  e�  s<  [� +  ,3       .    ,  s<  y  kl  y  kl  ��  s<  ��  s<  y +  ,4       .    ,  s<  e�  kl  e�  kl  y  s<  y  s<  e�      0    ,  c�  kl  [�  kl  [�  s<  c�  s<  c�  kl      1    ,  g�  g�  W�  g�  W�  w$  g�  w$  g�  g� +  ,5       .    ,  S�  [�  L,  [�  L,  e�  S�  e�  S�  [� +  ,6       .    ,  S�  y  L,  y  L,  ��  S�  ��  S�  y +  ,7       .    ,  S�  e�  L,  e�  L,  y  S�  y  S�  e�      0    ,  D\  kl  <�  kl  <�  s<  D\  s<  D\  kl      1    ,  HD  g�  8�  g�  8�  w$  HD  w$  HD  g� +  ,8       .    ,  4�  [�  ,�  [�  ,�  e�  4�  e�  4�  [� +  ,9       .    ,  4�  y  ,�  y  ,�  ��  4�  ��  4�  y +  ,10      .    ,  4�  e�  ,�  e�  ,�  y  4�  y  4�  e�      0    ,  %  kl  L  kl  L  s<  %  s<  %  kl      1    ,  )  g�  d  g�  d  w$  )  w$  )  g� +  ,11      +    ,  ��  e�  p  e�  p  y  ��  y  ��  e�      )    ,  �(  N       N       ��  �(  ��  �(  N  +  ,13      -    ,  ��  ]�  �  ]�  �  ��  ��  ��  ��  ]�      +    ,  ,�  e�  p  e�  p  y  ,�  y  ,�  e� +  ,12   
  via    6�  �   
  via    ��  �   
  via    Y�  �      3    ,  ,�  �P  @t  �P  @t  ��  ,�  ��  ,�  �P      3    ,  y  �P  ��  �P  ��  ��  y  ��  y  �P      3    ,  P  �P  c�  �P  c�  ��  P  ��  P  �P      1    ,     ��  �( ��  �( ��     ��     ��      1    ,          �(      �(  '      '              1    ,          �(      �(  '      '              1    ,     ��  �( ��  �( ��     ��     ��      �    ,          �(      �( ��     ��           	   1      � $  ��  ��  �� �  { �  { 4      1    ,  N   �D  ]�  �D  ]�  ��  N   ��  N   �D   	   1      � $  ~�  �P  ~�  ��  a�  ��  a�  w$   	   1      �   X &�  X  kl   	   1      �   a�  �$  !4  �$      1    ,  .�  �D  >�  �D  >�  ��  .�  ��  .�  �D      1    ,  a�  �T  qH  �T  qH  ��  a�  ��  a�  �T      1    ,  :� Y�  HD Y�  HD m<  :� m<  :� Y�      1    ,  :� m<  J8 m<  J8 ��  :� ��  :� m<      1    ,  :�  S�  FP  S�  FP  g�  :�  g�  :�  S�      1    ,  w$  '  ��  '  ��  S�  w$  S�  w$  '      1    ,  y  S�  ��  S�  ��  g�  y  g�  y  S�      1    ,  8�  '  HD  '  HD  S�  8�  S�  8�  '      )    ,      '  �(  '  �(  ��      ��      '      )    ,          �(      �(  *�      *�              *    ,     �  �( �  �( ��     ��     �      *    ,     ��  �( ��  �( ��     ��     ��   	   .      �   0� |  0�  ��      .    ,  _�  �`  s<  �`  s<  ��  _�  ��  _�  �`   	   .      �   U� |  P |  P  ��      .    ,  ,�  �P  @t  �P  @t  ��  ,�  ��  ,�  �P   	   .      �   oT  �`  oT  ��   	   .      �   ix |  ix  ��      .    ,  L,  �P  _�  �P  _�  ��  L,  ��  L,  �P      /    ,  2�  �,  :�  �,  :�  ��  2�  ��  2�  �,      /    ,  e�  �<  m`  �<  m`  �  e�  �  e�  �<      /    ,  R  �,  Y�  �,  Y�  ��  R  ��  R  �,              P  � GND  +  ,1               P �8 VDD  +  ,1               6�  � A1 +  ,1               ��  � Y  +  ,1               Y�  � A0 +  ,1       -    ,  0� cx  S� cx  S� ��  0� ��  0� cx      -    ,  � ��  �� ��  �� ��  � ��  � ��      ,    ,  .�  *�  R  *�  R  ]�  .�  ]�  .�  *�      ,    ,  m`  *�  ��  *�  ��  ]�  m`  ]�  m`  *�      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      +    ,  p ��  �� ��  �� �   p �   p ��      +    ,  6�  #(  J8  #(  J8  U�  6�  U�  6�  #(      +    ,  8� [�  J8 [�  J8 kH  8� kH  8� [�      +    ,  8� kH  L, kH  L, ��  8� ��  8� kH      +    ,  w$  U�  ��  U�  ��  e�  w$  e�  w$  U�      +    ,  8�  U�  HD  U�  HD  e�  8�  e�  8�  U�      +    ,  u0  #(  ��  #(  ��  U�  u0  U�  u0  #(      +    ,  p  �  ��  �  ��  #(  p  #(  p  �      0    ,  L �t  % �t  % �D  L �D  L �t      0    ,  <�  HD  D\  HD  D\  P  <�  P  <�  HD      0    ,  L  |  %  |  %  L  L  L  L  |      0    ,  4�  |  <�  |  <�  L  4�  L  4�  |      0    ,  L,  |  S�  |  S�  L  L,  L  L,  |      0    ,  c�  |  kl  |  kl  L  c�  L  c�  |      0    ,  {  HD  ��  HD  ��  P  {  P  {  HD      0    ,  <�  0�  D\  0�  D\  8�  <�  8�  <�  0�      0    ,  { �t  �� �t  �� �D  { �D  { �t      0    ,  c� �t  kl �t  kl �D  c� �D  c� �t      0    ,  L, �t  S� �t  S� �D  L, �D  L, �t      0    ,  4� �t  <� �t  <� �D  4� �D  4� �t      0    ,  >� ��  FP ��  FP �d  >� �d  >� ��      0    ,  >� q$  FP q$  FP x�  >� x�  >� q$      0    ,  >� �  FP �  FP ��  >� ��  >� �      0    ,  {  0�  ��  0�  ��  8�  {  8�  {  0�      0    ,  {  |  ��  |  ��  L  {  L  {  |              P  � GND               P �8 VDD               6�  � A1              ��  � Y               Y�  � A0     �     -� 	   0 9 
oai21     +    ,  �� 	�  s< 	�  s< z�  �� z�  �� 	� +  ,2       0    ,  �� |  { |  { L  �� L  �� |      0    ,  �� &�  { &�  { .�  �� .�  �� &�      0    ,  �� >\  { >\  { F,  �� F,  �� >\      0    ,  �� U�  { U�  { ]�  �� ]�  �� U�      0    ,  �� m<  { m<  { u  �� u  �� m<      1    ,  �� �  w$ �  w$ x�  �� x�  �� � +  ,1       .    ,  s<  ��  kl  ��  kl 	�  s< 	�  s<  �� +  ,3       .    ,  s< z�  kl z�  kl ��  s< ��  s< z� +  ,4       .    ,  s< 	�  kl 	�  kl z�  s< z�  s< 	�      .    ,  [�  ��  S�  ��  S� 	�  [� 	�  [�  �� +  ,5       .    ,  [� z�  S� z�  S� ��  [� ��  [� z� +  ,6       .    ,  [� 	�  S� 	�  S� z�  [� z�  [� 	�      0    ,  L, |  D\ |  D\ L  L, L  L, |      0    ,  L, &�  D\ &�  D\ .�  L, .�  L, &�      0    ,  L, >\  D\ >\  D\ F,  L, F,  L, >\      0    ,  L, U�  D\ U�  D\ ]�  L, ]�  L, U�      0    ,  L, m<  D\ m<  D\ u  L, u  L, m<      1    ,  P �  @t �  @t x�  P x�  P � +  ,7       .    ,  :�  ��  2�  ��  2� 	�  :� 	�  :�  �� +  ,8       .    ,  :� D8  2� D8  2� M�  :� M�  :� D8 +  ,9       .    ,  :� 	�  2� 	�  2� D8  :� D8  :� 	�      0    ,  *�   #(   #( &�  *� &�  *�       0    ,  *� 6�  #( 6�  #( >\  *� >\  *� 6�      1    ,  .� 4  @ 4  @ BD  .� BD  .� 4 +  ,10      +    L  #( 	�  #( @  L @  L D8  >� D8  >� z�  �� z�  �� 	�  #( 	�      *    L  �  �0  � �  � �  � [�  ' [�  ' �X  �( �X  �(  �0  �  �0 +  ,12      ,    L  X �  X p  | p  | L  6� L  6� ��  �� ��  �� �  X �      +    <  #( 	�  #( @  L @  L D8  2� D8  2� 	�  #( 	� +  ,11      +    ,  p  a�  ,�  a�  ,�  ��  p  ��  p  a� +  ,2       0    ,  L  g�  %  g�  %  oT  L  oT  L  g�      0    ,  L  ~�  %  ~�  %  ��  L  ��  L  ~�      1    ,  d  c�  )  c�  )  ��  d  ��  d  c� +  ,1       .    ,  ,�  W�  4�  W�  4�  a�  ,�  a�  ,�  W� +  ,3       .    ,  ,�  ��  4�  ��  4�  �d  ,�  �d  ,�  �� +  ,4       .    ,  ,�  a�  4�  a�  4�  ��  ,�  ��  ,�  a�      0    ,  <�  g�  D\  g�  D\  oT  <�  oT  <�  g�      0    ,  <�  ~�  D\  ~�  D\  ��  <�  ��  <�  ~�      1    ,  8�  c�  HD  c�  HD  ��  8�  ��  8�  c� +  ,5       .    ,  L,  W�  S�  W�  S�  a�  L,  a�  L,  W� +  ,6       .    ,  L,  ��  S�  ��  S�  �d  L,  �d  L,  �� +  ,7       .    ,  L,  a�  S�  a�  S�  ��  L,  ��  L,  a�      0    ,  [�  g�  c�  g�  c�  oT  [�  oT  [�  g�      0    ,  [�  ~�  c�  ~�  c�  ��  [�  ��  [�  ~�      1    ,  W�  c�  g�  c�  g�  ��  W�  ��  W�  c� +  ,8       .    ,  kl  W�  s<  W�  s<  a�  kl  a�  kl  W� +  ,9       .    ,  kl  ��  s<  ��  s<  �d  kl  �d  kl  �� +  ,10      .    ,  kl  a�  s<  a�  s<  ��  kl  ��  kl  a�      0    ,  {  g�  ��  g�  ��  oT  {  oT  {  g�      0    ,  {  ~�  ��  ~�  ��  ��  {  ��  {  ~�      1    ,  w$  c�  ��  c�  ��  ��  w$  ��  w$  c� +  ,11      +    ,  p  a�  ��  a�  ��  ��  p  ��  p  a�      )    ,      J8  �(  J8  �(  �      �      J8 +  ,13      -    ,  �  Y�  ��  Y�  ��  �p  �  �p  �  Y�      +    ,  s<  a�  ��  a�  ��  ��  s<  ��  s<  a� +  ,12   
  via    <�  �   
  via    _�  �   
  via    ��  �   
  via    d  �      3    ,  U�  �P  ix  �P  ix  ��  U�  ��  U�  �P      3    ,  y  �P  ��  �P  ��  ��  y  ��  y  �P      3    ,  2�  �P  FP  �P  FP  ��  2�  ��  2�  �P      3    ,  �  �P  #(  �P  #(  ��  �  ��  �  �P      1    ,          �(      �(  '      '              1    ,     ��  �( ��  �( ��     ��     ��      �    ,          �(      �( ��     ��              .    ,  y  �P  ��  �P  ��  ��  y  ��  y  �P      .    ,  2�  �P  FP  �P  FP  ��  2�  ��  2�  �P      .    ,  �  �P  #(  �P  #(  ��  �  ��  �  �P   	   .      �   :�  ��  @  ��  @  ��   	   .      �   kl  ��  }   ��  }   ��   	   .      � $  Bh  ��  Bh  �l  W�  �l  W�  ��   	   .      �   kl  �L  }   �L  }   �P   	   .      �   4�  �L  @  �L  @  �P   	   .      � $  Bh  �P  Bh  ��  P  ��  P  �d      /    ,  8�  �,  @t  �,  @t  ��  8�  ��  8�  �,      /    ,  ~�  �,  ��  �,  ��  ��  ~�  ��  ~�  �,      /    ,  |  �,  L  �,  L  ��  |  ��  |  �,      )    ,          �(      �(  �      �              *    ,      �0  �(  �0  �( ��     ��      �0      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      ,    ,  �  *�  2�  *�  2�  Y�  �  Y�  �  *�      -    ,  � ��  �� ��  �� ��  � ��  � ��      -    ,  m` ��  �� ��  �� ��  m` ��  m` ��      -    <  | L  6� L  6� ��  8� ��  8� ��  | ��  | L      1    ,  {  �D  ��  �D  ��  ��  {  ��  {  �D   	   1      �   _�  ��  _�  �P      1    ,  4�  �D  D\  �D  D\  ��  4�  ��  4�  �D      1    ,  d  R  '  R  '  c�  d  c�  d  R      1    ,  w$ �p  �� �p  �� ��  w$ ��  w$ �p   	   1      � $  @t  c�  @t  J8  ~�  J8  ~�  c�   	   1      � $  _�  ��  _�  �$  HD  �$  HD �      1    ,  �  �D  !4  �D  !4  ��  �  ��  �  �D      1    ,  d  '  )  '  )  R  d  R  d  '      1    ,  y x�  �� x�  �� �p  y �p  y x�      1    ,  @ BD  ,� BD  ,� U�  @ U�  @ BD      1    ,  @ U�  .� U�  .� ��  @ ��  @ U�      +    ,  p ��  �� ��  �� �   p �   p ��      +    ,  p  �  ��  �  ��  #(  p  #(  p  �      +    ,  p  S�  )  S�  )  a�  p  a�  p  S�      +    ,  p  #(  *�  #(  *�  S�  p  S�  p  #(      +    ,  w$ z�  �� z�  �� �|  w$ �|  w$ z�      +    ,  u0 �|  �� �|  �� ��  u0 ��  u0 �|      +    ,  L D8  .� D8  .� S�  L S�  L D8      +    ,  L S�  0� S�  0� ��  L ��  L S�      0    ,  4� �t  <� �t  <� �D  4� �D  4� �t      0    ,  L, �t  S� �t  S� �D  L, �D  L, �t      0    ,  { �t  �� �t  �� �D  { �D  { �t      0    ,  c� �t  kl �t  kl �D  c� �D  c� �t      0    ,  L �t  % �t  % �D  L �D  L �t      0    ,  c�  |  kl  |  kl  L  c�  L  c�  |      0    ,  L  |  %  |  %  L  L  L  L  |      0    ,  4�  |  <�  |  <�  L  4�  L  4�  |      0    ,  L,  |  S�  |  S�  L  L,  L  L,  |      0    ,  {  |  ��  |  ��  L  {  L  {  |      0    ,  L  FP  %  FP  %  N   L  N   L  FP      0    ,  L  .�  %  .�  %  6�  L  6�  L  .�      0    ,  { �X  �� �X  �� �(  { �(  { �X      0    ,  #( q$  *� q$  *� x�  #( x�  #( q$      0    ,  #( ��  *� ��  *� �d  #( �d  #( ��      0    ,  #( �  *� �  *� ��  #( ��  #( �      0    ,  #( Y�  *� Y�  *� a�  #( a�  #( Y�              P  � GND  +  ,1               P �8 VDD  +  ,1               ��  � A0 +  ,1               <�  � A1 +  ,1               _�  � Y  +  ,1               d  � B0 +  ,1               P  � GND               P �8 VDD               ��  � A0              <�  � A1              _�  � Y               d  � B0     �   
  	� 	   /  
aoi22     0    ,  �   �L   �L &�  � &�  �       0    ,  � 6�  �L 6�  �L >\  � >\  � 6�      0    ,  � M�  �L M�  �L U�  � U�  � M�      1    ,  � 4  �d 4  �d Y�  � Y�  � 4 +  ,1       .    ,  �| |  �� |  �� @  �| @  �| | +  ,3       .    ,  �| [�  �� [�  �� el  �| el  �| [� +  ,4       .    ,  �| @  �� @  �� [�  �| [�  �| @      0    ,  ��   {   { &�  �� &�  ��       0    ,  �� 6�  { 6�  { >\  �� >\  �� 6�      0    ,  �� M�  { M�  { U�  �� U�  �� M�      1    ,  �� 4  w$ 4  w$ Y�  �� Y�  �� 4 +  ,5       .    ,  s< |  kl |  kl @  s< @  s< | +  ,6       .    ,  s< [�  kl [�  kl el  s< el  s< [� +  ,7       .    ,  s< @  kl @  kl [�  s< [�  s< @      0    ,  c�   [�   [� &�  c� &�  c�       0    ,  c� 6�  [� 6�  [� >\  c� >\  c� 6�      0    ,  c� M�  [� M�  [� U�  c� U�  c� M�      1    ,  g� 4  W� 4  W� Y�  g� Y�  g� 4 +  ,8       .    ,  S� |  L, |  L, @  S� @  S� | +  ,9       .    ,  S� [�  L, [�  L, el  S� el  S� [� +  ,10      .    ,  S� @  L, @  L, [�  S� [�  S� @      0    ,  D\   <�   <� &�  D\ &�  D\       0    ,  D\ 6�  <� 6�  <� >\  D\ >\  D\ 6�      0    ,  D\ M�  <� M�  <� U�  D\ U�  D\ M�      1    ,  HD 4  8� 4  8� Y�  HD Y�  HD 4 +  ,11      .    ,  4� |  ,� |  ,� @  4� @  4� | +  ,12      .    ,  4� [�  ,� [�  ,� el  4� el  4� [� +  ,13      .    ,  4� @  ,� @  ,� [�  4� [�  4� @      0    ,  %   L   L &�  % &�  %       0    ,  % 6�  L 6�  L >\  % >\  % 6�      0    ,  % M�  L M�  L U�  % U�  % M�      1    ,  ) 4  d 4  d Y�  ) Y�  ) 4 +  ,14      +    ,  �� @  p @  p [�  �� [�  �� @      +    ,  �� @  �| @  �| [�  �� [�  �� @ +  ,2       *    ,  �h �     �     s  �h s  �h � +  ,16      ,    ,  �� p  � p  � cx  �� cx  �� p      +    ,  ,� @  p @  p [�  ,� [�  ,� @ +  ,15      +    ,  �(  e�  ��  e�  ��  ��  �(  ��  �(  e� +  ,2       0    ,  �L  kl  �|  kl  �|  s<  �L  s<  �L  kl      0    ,  �L  ��  �|  ��  �|  ��  �L  ��  �L  ��      1    ,  �4  g�  ��  g�  ��  ��  �4  ��  �4  g� +  ,1       .    ,  ��  [�  ��  [�  ��  e�  ��  e�  ��  [� +  ,3       .    ,  ��  ��  ��  ��  ��  �L  ��  �L  ��  �� +  ,4       .    ,  ��  e�  ��  e�  ��  ��  ��  ��  ��  e�      .    ,  s<  [�  kl  [�  kl  e�  s<  e�  s<  [� +  ,5       .    ,  s<  ��  kl  ��  kl  �L  s<  �L  s<  �� +  ,6       .    ,  s<  e�  kl  e�  kl  ��  s<  ��  s<  e�      0    ,  c�  kl  [�  kl  [�  s<  c�  s<  c�  kl      0    ,  c�  ��  [�  ��  [�  ��  c�  ��  c�  ��      1    ,  g�  g�  W�  g�  W�  ��  g�  ��  g�  g� +  ,7       .    ,  S�  [�  L,  [�  L,  e�  S�  e�  S�  [� +  ,8       .    ,  S�  ��  L,  ��  L,  �L  S�  �L  S�  �� +  ,9       .    ,  S�  e�  L,  e�  L,  ��  S�  ��  S�  e�      .    ,  <�  [�  4�  [�  4�  e�  <�  e�  <�  [� +  ,10      .    ,  <�  ��  4�  ��  4�  �L  <�  �L  <�  �� +  ,11      .    ,  <�  e�  4�  e�  4�  ��  <�  ��  <�  e�      0    ,  ,�  kl  %  kl  %  s<  ,�  s<  ,�  kl      0    ,  ,�  ��  %  ��  %  ��  ,�  ��  ,�  ��      1    ,  0�  g�  !4  g�  !4  ��  0�  ��  0�  g� +  ,12      +    ,  �(  e�  @  e�  @  ��  �(  ��  �(  e�      )    ,  ��  N   �  N   �  ��  ��  ��  ��  N  +  ,14      -    ,  ��  ]�  p  ]�  p  �X  ��  �X  ��  ]�      +    ,  4�  e�  @  e�  @  ��  4�  ��  4�  e� +  ,13   
  via  �  B�         d  �   
  via  �  B�         <�  �   
  via  �  B�         _�  �   
  via  �  B�         ��  �   
  via  �  B�         �  �      1    ,     ��  �h ��  �h ��     ��     ��      1    ,          �h      �h  '      '              1    ,     ��  �h ��  �h ��     ��     ��      1    ,          �h      �h  '      '              3    ,  �  �P  #(  �P  #(  ��  �  ��  �  �P      3    ,  2�  �P  FP  �P  FP  ��  2�  ��  2�  �P      3    ,  y  �P  ��  �P  ��  ��  y  ��  y  �P      3    ,  U�  �P  ix  �P  ix  ��  U�  ��  U�  �P      3    ,  �@  �P  ��  �P  ��  ��  �@  ��  �@  �P      /    ,  ~�  �,  ��  �,  ��  ��  ~�  ��  ~�  �,      /    ,  8�  �,  @t  �,  @t  ��  8�  ��  8�  �,      /    ,  [�  �,  c�  �,  c�  ��  [�  ��  [�  �,      /    ,  �  �,  ��  �,  ��  ��  �  ��  �  �,      )    ,          �h      �h  ��      ��              *    ,     �  �h �  �h ��     ��     �      ,    ,  �  �  ��  �  ��  *�  �  *�  �  �      ,    ,  ��  *�  ��  *�  ��  ]�  ��  ]�  ��  *�      ,    ,  p  *�  :�  *�  :�  ]�  p  ]�  p  *�      -    ,  � ��  �� ��  �� ��  � ��  � ��      -    ,  m` cx  �� cx  �� ��  m` ��  m` cx      +    ,  �  �  ��  �  ��  #(  �  #(  �  �      +    ,  � ��  �� ��  �� �   � �   � ��      +    ,  ��  U�  �(  U�  �(  e�  ��  e�  ��  U�      +    ,  ��  #(  �(  #(  �(  U�  ��  U�  ��  #(      +    ,  @  #(  2�  #(  2�  U�  @  U�  @  #(      +    ,  @  U�  0�  U�  0�  e�  @  e�  @  U�      +    ,  u0 kH  �� kH  �� ��  u0 ��  u0 kH      +    ,  w$ [�  �� [�  �� kH  w$ kH  w$ [�   	   1      � $  a� 4  a� �  �@ �  �@ 4   	   1      � $  >� 4  >�  ��  L  ��  L  ��   	   1      � $  ]� Y�  ]� s  #( s  #( Y�      1    ,  4�  �D  D\  �D  D\  ��  4�  ��  4�  �D      1    ,  �4  �D  ��  �D  ��  ��  �4  ��  �4  �D   	   1      � $  L  �P  L  ��  ]�  ��  ]�  ��      1    ,  {  �D  ��  �D  ��  ��  {  ��  {  �D      1    ,  W�  �D  g�  �D  g�  ��  W�  ��  W�  �D      1    ,  ��  S�  �4  S�  �4  g�  ��  g�  ��  S�      1    ,  ��  '  �4  '  �4  S�  ��  S�  ��  '      1    ,  !4  '  0�  '  0�  S�  !4  S�  !4  '      1    ,  !4  S�  .�  S�  .�  g�  !4  g�  !4  S�      1    ,  y Y�  �� Y�  �� m<  y m<  y Y�      1    ,  w$ m<  �� m<  �� ��  w$ ��  w$ m<      0    ,  ,�  |  4�  |  4�  L  ,�  L  ,�  |      0    ,  D\  |  L,  |  L,  L  D\  L  D\  |      0    ,  [�  |  c�  |  c�  L  [�  L  [�  |      0    ,  s<  |  {  |  {  L  s<  L  s<  |      0    ,  ��  |  �|  |  �|  L  ��  L  ��  |      0    ,  |  |  L  |  L  L  |  L  |  |      0    ,  �  |  ��  |  ��  L  �  L  �  |      0    ,  | �t  L �t  L �D  | �D  | �t      0    ,  ,� �t  4� �t  4� �D  ,� �D  ,� �t      0    ,  D\ �t  L, �t  L, �D  D\ �D  D\ �t      0    ,  [� �t  c� �t  c� �D  [� �D  [� �t      0    ,  s< �t  { �t  { �D  s< �D  s< �t      0    ,  �� �t  �| �t  �| �D  �� �D  �� �t      0    ,  � �t  �� �t  �� �D  � �D  � �t      0    ,  �|  HD  �L  HD  �L  P  �|  P  �|  HD      0    ,  �|  0�  �L  0�  �L  8�  �|  8�  �|  0�      0    ,  %  0�  ,�  0�  ,�  8�  %  8�  %  0�      0    ,  %  HD  ,�  HD  ,�  P  %  P  %  HD      0    ,  { q$  �� q$  �� x�  { x�  { q$      0    ,  { ��  �� ��  �� �d  { �d  { ��      0    ,  { �  �� �  �� ��  { ��  { �      .    ,  y  �P  ��  �P  ��  ��  y  ��  y  �P      .    ,  �@  �P  ��  �P  ��  ��  �@  ��  �@  �P      .    ,  U�  �P  ix  �P  ix  ��  U�  ��  U�  �P      .    ,  2�  �P  FP  �P  FP  ��  2�  ��  2�  �P   	   .      �   8�  �L  8�  �P   	   .      � $  P |  P  �x  Y�  �x  Y�  ��   	   .      � $  �(  ��  �(  �   ��  �   �� |   	   .      � $  0� |  0�  �x  6�  �x  6�  ��   	   .      � $  oT |  oT  �x  }   �x  }   ��   	   .      � $  }   �P  }   ��  oT  ��  oT  �L   	   .      �   ��  �L  �(  �L  �(  �P   	   .      �   Y�  �P  Y�  �4  L,  �4              _�  � GND  +  ,1               _� �8 VDD  +  ,1               ��  � A0 +  ,1               _�  � B0 +  ,1               <�  � B1 +  ,1               �  � A1 +  ,1               d  � Y  +  ,1       �    ,          �h      �h ��     ��                      _�  � GND               _� �8 VDD               ��  � A0              _�  � B0              <�  � B1              �  � A1              d  � Y      �      � 	   1 . 
xnor2     +    ,  ި  Y�  �,  Y�  �,  ��  ި  ��  ި  Y� +  ,2       0    ,  ��  _�  ��  _�  ��  g�  ��  g�  ��  _�      0    ,  ��  w$  ��  w$  ��  ~�  ��  ~�  ��  w$      1    ,  ܴ  [�  �  [�  �  ��  ܴ  ��  ܴ  [� +  ,1       .    ,  �,  P  �\  P  �\  Y�  �,  Y�  �,  P +  ,3       .    ,  �,  ��  �\  ��  �\  ��  �,  ��  �,  �� +  ,4       .    ,  �,  Y�  �\  Y�  �\  ��  �,  ��  �,  Y�      0    ,  ��  _�  ��  _�  ��  g�  ��  g�  ��  _�      0    ,  ��  w$  ��  w$  ��  ~�  ��  ~�  ��  w$      1    ,  �t  [�  ��  [�  ��  ��  �t  ��  �t  [� +  ,5       .    ,  ��  P  �  P  �  Y�  ��  Y�  ��  P +  ,6       .    ,  ��  ��  �  ��  �  ��  ��  ��  ��  �� +  ,7       .    ,  ��  Y�  �  Y�  �  ��  ��  ��  ��  Y�      0    ,  �L  _�  �|  _�  �|  g�  �L  g�  �L  _�      0    ,  �L  w$  �|  w$  �|  ~�  �L  ~�  �L  w$      1    ,  �4  [�  ��  [�  ��  ��  �4  ��  �4  [� +  ,8       .    ,  ��  P  ��  P  ��  Y�  ��  Y�  ��  P +  ,9       .    ,  ��  ��  ��  ��  ��  ��  ��  ��  ��  �� +  ,10      .    ,  ��  Y�  ��  Y�  ��  ��  ��  ��  ��  Y�      0    ,  {  _�  s<  _�  s<  g�  {  g�  {  _�      0    ,  {  w$  s<  w$  s<  ~�  {  ~�  {  w$      1    ,  ~�  [�  oT  [�  oT  ��  ~�  ��  ~�  [� +  ,11      +    ,  ި  Y�  m`  Y�  m`  ��  ި  ��  ި  Y�      )    ,  �  Bh  U�  Bh  U�  �@  �  �@  �  Bh +  ,13      -    ,  �x  R  e�  R  e�  ��  �x  ��  �x  R      +    ,  ��  Y�  m`  Y�  m`  ��  ��  ��  ��  Y� +  ,12      +    ,  a�  Y�  L,  Y�  L,  ��  a�  ��  a�  Y� +  ,2       0    ,  [�  _�  S�  _�  S�  g�  [�  g�  [�  _�      0    ,  [�  w$  S�  w$  S�  ~�  [�  ~�  [�  w$      1    ,  _�  [�  P  [�  P  ��  _�  ��  _�  [� +  ,1       .    ,  L,  P  D\  P  D\  Y�  L,  Y�  L,  P +  ,3       .    ,  L,  ��  D\  ��  D\  ��  L,  ��  L,  �� +  ,4       .    ,  L,  Y�  D\  Y�  D\  ��  L,  ��  L,  Y�      .    ,  4�  P  ,�  P  ,�  Y�  4�  Y�  4�  P +  ,5       .    ,  4�  ��  ,�  ��  ,�  ��  4�  ��  4�  �� +  ,6       .    ,  4�  Y�  ,�  Y�  ,�  ��  4�  ��  4�  Y�      0    ,  %  _�  L  _�  L  g�  %  g�  %  _�      0    ,  %  w$  L  w$  L  ~�  %  ~�  %  w$      1    ,  )  [�  d  [�  d  ��  )  ��  )  [� +  ,7       +    ,  a�  Y�  p  Y�  p  ��  a�  ��  a�  Y�      )    ,  y  Bh      Bh      �@  y  �@  y  Bh +  ,9       -    ,  ix  R  �  R  �  ��  ix  ��  ix  R      +    ,  ,�  Y�  p  Y�  p  ��  ,�  ��  ,�  Y� +  ,8       0    ,  8� �  @t �  @t �  8� �  8� �      0    ,  8� (  @t (  @t $�  8� $�  8� (      0    ,  8� 4�  @t 4�  @t <h  8� <h  8� 4�      1    ,  4� �  D\ �  D\ @P  4� @P  4� � +  ,1       .    ,  HD  �  P  �  P  ��  HD  ��  HD  � +  ,3       .    ,  HD BD  P BD  P L  HD L  HD BD +  ,4       .    ,  HD  ��  P  ��  P BD  HD BD  HD  ��      0    ,  W� �  _� �  _� �  W� �  W� �      0    ,  W� (  _� (  _� $�  W� $�  W� (      0    ,  W� 4�  _� 4�  _� <h  W� <h  W� 4�      1    ,  S� �  c� �  c� @P  S� @P  S� � +  ,5       .    ,  g�  �  oT  �  oT  ��  g�  ��  g�  � +  ,6       .    ,  g� BD  oT BD  oT L  g� L  g� BD +  ,7       .    ,  g�  ��  oT  ��  oT BD  g� BD  g�  ��      0    ,  y p  �� p  �� @  y @  y p      0    ,  y (�  �� (�  �� 0�  y 0�  y (�      0    ,  y @P  �� @P  �� H   y H   y @P      0    ,  y W�  �� W�  �� _�  y _�  y W�      0    ,  y o0  �� o0  �� w   y w   y o0      1    ,  u0 �  �� �  �� z�  u0 z�  u0 � +  ,8       .    ,  ��  �  ��  �  ��  ��  ��  ��  ��  � +  ,9       .    ,  �� |�  �� |�  �� ��  �� ��  �� |� +  ,10      .    ,  ��  ��  ��  ��  �� |�  �� |�  ��  ��      .    ,  �(  �  ��  �  ��  ��  �(  ��  �(  � +  ,11      .    ,  �( |�  �� |�  �� ��  �( ��  �( |� +  ,12      .    ,  �(  ��  ��  ��  �� |�  �( |�  �(  ��      0    ,  �� �  �� �  �� �  �� �  �� �      0    ,  �� (  �� (  �� $�  �� $�  �� (      0    ,  �� 4�  �� 4�  �� <h  �� <h  �� 4�      0    ,  �� L  �� L  �� S�  �� S�  �� L      0    ,  �� cx  �� cx  �� kH  �� kH  �� cx      1    ,  �� �  �� �  �� o0  �� o0  �� � +  ,13      .    ,  �\  �  �,  �  �,  ��  �\  ��  �\  � +  ,14      .    ,  �\ BD  �, BD  �, L  �\ L  �\ BD +  ,15      .    ,  �\  ��  �,  ��  �, BD  �\ BD  �\  ��      0    ,  �� �  �� �  �� �  �� �  �� �      0    ,  �� (  �� (  �� $�  �� $�  �� (      0    ,  �� 4�  �� 4�  �� <h  �� <h  �� 4�      1    ,  � �  ܴ �  ܴ @P  � @P  � � +  ,16      +    \  ި  ��  ި BD  �t BD  �t q$  �� q$  �� |�  s< |�  s< BD  2� BD  2�  ��  ި  ��      *    \  �  �l  � Y�  �� Y�  �� ��  � ��  � �L  [� �L  [� Y�  X Y�  X  �l  �  �l +  ,18      ,    \  �x  �  �x J  �D J  �D x�  �h x�  �h ��  kl ��  kl J  *� J  *�  �  �x  �      +    ,  2�  ��  HD  ��  HD BD  2� BD  2�  �� +  ,2       +    ,  �,  ��  ި  ��  ި BD  �, BD  �,  �� +  ,17   
  via    6�  �   
  via  �  B�         ��  �   
  via    ܴ  �      1    ,          �      �  '      '              1    ,     ��  � ��  � ��     ��     ��      3    ,  ,�  �P  @t  �P  @t  ��  ,�  ��  ,�  �P      3    ,  ��  �P  �X  �P  �X  ��  ��  ��  ��  �P      3    ,  ��  �P  �x  �P  �x  ��  ��  ��  ��  �P      �    ,          �      � ��     ��              )    ,          �      �  �@      �@              *    ,      �l  �  �l  � ��     ��      �l      ,    ,  �  �  �`  �  �`  *�  �  *�  �  �      ,    ,  FP  *�  ix  *�  ix  R  FP  R  FP  *�      ,    ,  �P  *�  �x  *�  �x  R  �P  R  �P  *�      0    ,  �t  |  �D  |  �D  L  �t  L  �t  |      0    ,  d  |  !4  |  !4  L  d  L  d  |      0    ,  0�  |  8�  |  8�  L  0�  L  0�  |      0    ,  HD  |  P  |  P  L  HD  L  HD  |      0    ,  _�  |  g�  |  g�  L  _�  L  _�  |      0    ,  w$  |  ~�  |  ~�  L  w$  L  w$  |      0    ,  ��  |  �d  |  �d  L  ��  L  ��  |      0    ,  �  |  ��  |  ��  L  �  L  �  |      0    ,  ��  |  ܴ  |  ܴ  L  ��  L  ��  |      0    ,  HD �t  P �t  P �D  HD �D  HD �t      0    ,  0� �t  8� �t  8� �D  0� �D  0� �t      0    ,  d �t  !4 �t  !4 �D  d �D  d �t      0    ,  _� �t  g� �t  g� �D  _� �D  _� �t      0    ,  w$ �t  ~� �t  ~� �D  w$ �D  w$ �t      0    ,  �� �t  �d �t  �d �D  �� �D  �� �t      0    ,  � �t  �� �t  �� �D  � �D  � �t      0    ,  �t �t  �D �t  �D �D  �t �D  �t �t      0    ,  �� �t  ܴ �t  ܴ �D  �� �D  �� �t      0    ,  S�  <�  [�  <�  [�  D\  S�  D\  S�  <�      0    ,  �� W�  �� W�  �� _�  �� _�  �� W�      0    ,  ��  <�  ��  <�  ��  D\  ��  D\  ��  <�      0    ,  8� o0  @t o0  @t w   8� w   8� o0      0    ,  8� ��  @t ��  @t �p  8� �p  8� ��      0    ,  8� �  @t �  @t ��  8� ��  8� �      0    ,  y �d  �� �d  �� �4  y �4  y �d      0    ,  �� o0  �� o0  �� w   �� w   �� o0      0    ,  �� ��  �� ��  �� �p  �� �p  �� ��      0    ,  �� �  �� �  �� ��  �� ��  �� �      0    ,  8� W�  @t W�  @t _�  8� _�  8� W�      +    ,  �  �  �  �  �  #(  �  #(  �  �      +    ,  � ��  � ��  � �   � �   � ��      +    ,  N   6�  a�  6�  a�  J8  N   J8  N   6�      +    ,  P  J8  a�  J8  a�  Y�  P  Y�  P  J8      +    ,  � BD  ި BD  ި Q�  � Q�  � BD      +    ,  s< ��  �� ��  �� �  s< �  s< ��      +    ,  �  J8  ި  J8  ި  Y�  �  Y�  �  J8      +    ,  �   #(  ި  #(  ި  J8  �   J8  �   #(      +    ,  s< |�  �� |�  �� ��  s< ��  s< |�      +    ,  2� Q�  FP Q�  FP ��  2� ��  2� Q�      +    ,  �  Q�  ި Q�  ި ��  �  ��  �  Q�      +    ,  2� BD  D\ BD  D\ Q�  2� Q�  2� BD   	   .      �   �  �  �  ��  �X  ��   	   .      �   0�  ��  0�  �P   	   .      �   ��  �|  D\  �|   	   .      � $  0�  P  0�  .�  �  .�  �  P   	   .      � $  ��  �  ��  �x  L,  �x  L,  �   	   .      �   ��  �d  ��  �    	   .      � $  � ��  � ��  kl ��  kl L   	   .      �   HD  �x  <�  �x  <�  ��      .    ,  ��  �P  �X  �P  �X  ��  ��  ��  ��  �P      .    ,  ,�  �P  @t  �P  @t  ��  ,�  ��  ,�  �P   	   .      �   �D  �  �D  ��      .    ,  ��  �  �8  �  �8  ��  ��  ��  ��  �      /    ,  2�  �,  :�  �,  :�  ��  2�  ��  2�  �,      /    ,  ��  �,  �|  �,  �|  ��  ��  ��  ��  �,      /    ,  ��  ��  �\  ��  �\  ��  ��  ��  ��  ��      -    ,  � ��  �` ��  �` ��  � ��  � ��      -    ,  kl ��  �� ��  �� ��  kl ��  kl ��      -    <  �h x�  �D x�  �D J  �x J  �x ��  �h ��  �h x�      -    ,  *� J  N  J  N  ��  *� ��  *� J      1    ,  u0 z�  �� z�  �� �|  u0 �|  u0 z�      1    ,  .�  �D  >�  �D  >�  ��  .�  ��  .�  �D      1    ,  P  8�  _�  8�  _�  HD  P  HD  P  8�      1    ,  P  '  _�  '  _�  8�  P  8�  P  '      1    ,  R  HD  _�  HD  _�  [�  R  [�  R  HD      1    ,  u0 �|  �� �|  �� �  u0 �  u0 �|      1    ,  � @P  ܴ @P  ܴ S�  � S�  � @P      1    ,  ��  �D  �d  �D  �d  ��  ��  ��  ��  �D      1    ,  � S�  ܴ S�  ܴ ��  � ��  � S�   	   1      �   [� �  [�  ��      1    ,  u0 �  �� �  �� ��  u0 ��  u0 �   	   1      �   ��  ��  !4  ��  !4  ��      1    ,  4� @P  Bh @P  Bh S�  4� S�  4� @P      1    ,  �  '  ܴ  '  ܴ  HD  �  HD  �  '      1    ,  �  HD  ܴ  HD  ܴ  [�  �  [�  �  HD   	   1      � $  ��  [�  ��  D\  w$  D\  w$  [�      1    ,  4� S�  D\ S�  D\ ��  4� ��  4� S�      1    ,  ��  ��  �D  ��  �D  ��  ��  ��  ��  ��   	   1      � $  �� �  ��  �T  ��  �T  ��  ��   	   1      � $  ��  �P  ��  �d  �d  �d  �d  ��              {  � GND  +  ,1               { �8 VDD  +  ,1               6�  � A0 +  ,1               ܴ  � Y  +  ,1               ��  � A1 +  ,1               {  � GND               { �8 VDD               6�  � A0              ܴ  � Y               ��  � A1     �    # 4�      
layout 
  
oai32   �@ #� +  
,ix3821   
  
buf02   �@ 
ɸ +  
,ix3714   
  
buf02  �  B�        �\ 
ɸ +  
,ix3716   
  
aoi21  �  B�        ^( tX +  
,ix3915   
  
aoi221  �@ � +  
,ix3474   
  
aoi221 �  B�        (( tX +  
,ix3442   
  
aoi221  
�@ � +  
,ix3506   
  
aoi221 �  B�        
�� tX +  
,ix3494   
  
aoi221  	G  � +  
,ix3526   
  
aoi221 �  B�        �h tX +  
,ix3410   
  
aoi221  �@ 
ɸ +  
,ix1684   
  
aoi221 �  B�        �h tX +  
,ix3430   
  
aoi221 �  B�        �h 
ɸ +  
,ix3462   
  ao22 �  B�        
�\ 
ɸ +  
,ix3547   
  ao22 �  B�        	�\ 
ɸ +  
,ix3491   
  ao22 �  B�        �� 
ɸ +  
,ix3905   
  ao22  $@ � +  
,ix3659   
  ao22 �  B�        �\ 
ɸ +  
,ix3603   
  
oai22  �  B�        �( /  +  
,ix3885   
  
oai22   �  /  +  
,ix3893   
  
oai22  �  B�        � Č +  
,ix3829   
  
oai22   y� �� +  
,ix3837   
  
oai22  �  B�        �(  X +  
,ix3845   
  
oai22   �@  X +  
,ix3853   
  
oai22  �  B�        �(  X +  
,ix3861   
  
oai22   K� "� +  
,ix3869   
  
oai22   E� l� +  
,ix3877   
  
oai22  �  B�        �� � +  
,ix3575   
  
oai22  �  B�        � tX +  
,ix3631   
  
oai22  �  B�        �� � +  
,ix3519   
  
oai22   �� tX +  
,ix3695   
  dffs_ni   )�  %$ +  ,fsm_inst_reg_state_0   
  or03  )#@ %$ +  ,ix13   
  
and02  �  B�        � l� +  
,ix3473   
  
and02  �  B�        � � +  
,ix3687   
  
and02  �  B�        -̜ #� +  ,ix19   
  dffr  *<� #� +  ,fsm_inst_reg_state_1   
  dffr �  B�        *!( #� +  ,fsm_inst_reg_state_2   
  dffr �  B�        (� %$ +  ,fsm_inst_reg_state_3   
  dffr �  B�        %�� %$ +  ,fsm_inst_reg_state_4   
  
nor02   �� "� +  
,ix3699   
  
nor02   #  tX +  
,ix3312   
  
nor02   Q� � +  
,ix3747   
  
nor02  �  B�        h 
ɸ +  
,ix3302   
  
nor02   � 
ɸ +  
,ix2466   
  
nor02  �  B�        )�( l� +  
,ix3154   
  
nor02   �� tX +  
,ix2076   
  
nor02   &s�  X +  
,ix3258   
  
nor02  �  B�        '� /  +  
,ix3262   
  
inv01  �  B�        	+�  X +  
,ix3632   
  
inv01  �  B�        (  X +  
,ix3564   
  
inv01   K�  X +  
,ix3628   
  
inv01   &� "� +  
,ix3556   
  
inv01    � l� +  
,ix3624   
  
inv01  �  B�        $h /  +  
,ix3548   
  
inv01  �  B�        $�� l� +  
,ix1517   
  
inv01  �  B�        r� "� +  
,ix3633   
  
inv01   8� l� +  
,ix3101   
  
inv01  �  B�        �( "� +  
,ix3406   
  
inv01   @ ! +  
,ix3642   
  
inv01   @ #� +  
,ix3803   
  
inv01  �  B�        � s4 +  
,ix3580   
  
inv01  �  B�        R( Č +  
,ix3636   
  
inv01  �  B�        �h "� +  
,ix3572   
  
inv01   
�  /  +  
,ix3620   
  
inv01  �  B�        4( tX +  
,ix3718   
  
inv01  �  B�        �( tX +  
,ix3720   
  
inv01   �  � +  
,ix3308   
  
inv01  �  B�         � � +  
,ix1341   
  
inv01   N@ � +  
,ix2937   
  
inv01     � +  
,ix3689   
  
inv01   6@ l� +  
,ix3738   
  
inv01   
!� l� +  
,ix3740   
  
inv01   �@ � +  
,ix1393   
  
inv01  �  B�        �( tX +  
,ix2989   
  
inv01  �  B�        �( tX +  
,ix3734   
  
inv01   S  tX +  
,ix3736   
  
inv01  �  B�        �( 
ɸ +  
,ix1289   
  
inv01   
`@ � +  
,ix2885   
  
inv01  �  B�        �h l� +  
,ix3041   
  
inv01  �  B�        �� "� +  
,ix3521   
  
inv01   	� "� +  
,ix3577   
  
inv01  �  B�        :( tX +  
,ix3679   
  
inv01  �  B�        � tX +  
,ix3467   
  
inv01  �  B�         � tX +  
,ix3685   
  
inv01   �@ � +  
,ix3314   
  
inv01  �  B�        /h tX +  
,ix1445   
  
inv01   
�� 8� +  
,ix3034   
  
inv01  �  B�        "�� �� +  
,ix2876   
  
inv01  �  B�         �� Č +  
,ix3046   
  
inv01   ƀ �T +  
,ix2868   
  
inv01   t� �T +  
,ix3040   
  
inv01   �@ �T +  
,ix1167   
  
inv01   Z@ �T +  
,ix3728   
  
inv01   M   +  
,ix997    
  
inv01   �� 8� +  
,ix991    
  
inv01  �  B�        �( s4 +  
,ix2858   
  
inv01   �� #� +  
,ix2566   
  
inv01   ؀ %$ +  
,ix2742   
  
inv01  �  B�        � 8� +  
,ix545    
  
inv01   *@ �d +  
,ix3726   
  
inv01   �  #� +  
,ix375    
  
inv01   �� ! +  
,ix369    
  
inv01    Y@ %$ +  
,ix2576   
  
inv01   !�@ %$ +  
,ix2748   
  
inv01  �  B�        )� ! +  
,ix2582   
  
inv01  �  B�        &�� ! +  
,ix2754   
  
inv01   H@ /  +  
,ix3730   
  
inv01   ~@ �� +  
,ix1959   
  
inv01   � Č +  
,ix1953   
  
inv01  �  B�        h �T +  
,ix2204   
  
inv01   �   +  
,ix2446   
  
inv01   H@ �� +  
,ix2214   
  
inv01   /  �T +  
,ix2424   
  
inv01  �  B�        Ѩ �� +  
,ix2222   
  
inv01  �  B�        �h /  +  
,ix2402   
  
inv01   �@ /  +  
,ix2129   
  
inv01  �  B�        ר 
ɸ +  
,ix1800   
  
inv01  �  B�        Z� /  +  
,ix1984   
  
inv01   �� Č +  
,ix1792   
  
inv01  �  B�        �� �� +  
,ix1978   
  
inv01   �� �T +  
,ix1782   
  
inv01   �� Č +  
,ix1972   
  
inv01   
�� l� +  
,ix2751   
  
inv01   	G  /  +  
,ix3732   
  
inv01  �  B�        �( �� +  
,ix2575   
  
inv01   Q� Č +  
,ix2581   
  
inv01  �  B�        *~� v� +  
,ix679    
  
inv01   �� /  +  
,ix1711   
  
inv01  �  B�        -�( 8� +  
,ix2492   
  
inv01  �  B�        .�( �d +  
,ix2494   
  
inv01  �  B�        �( s4 +  
,ix2792   
  
inv01  �  B�        �� s4 +  
,ix2500   
  
inv01  �  B�        �( ! +  
,ix2798   
  
inv01  �  B�        Ѩ ! +  
,ix2506   
  
inv01   ,O� �T +  ,ix57   
  
inv01   +�@ v� +  
,ix749    
  
inv01   %y�  +  
,ix1710   
  
inv01     8� +  
,ix1716   
  
inv01   Q� s4 +  
,ix1722   
  
inv01  �  B�        U� v� +  
,ix1641   
  
inv01  �  B�        #+� 
ɸ +  
,ix2427   
  
inv01  �  B�        "�( v� +  
,ix1876   
  
inv01   �� �T +  
,ix2140   
  
inv01  �  B�        [� 8� +  
,ix1908   
  
inv01  �  B�        h ! +  
,ix2146   
  
inv01  �  B�        �h %$ +  
,ix1938   
  
inv01  �  B�        	h %$ +  
,ix2152   
  
inv01  �  B�        -ʨ  +  
,ix127    
  
inv01  �  B�         |h v� +  
,ix1875   
  
inv01  �  B�        -l� �� +  
,ix2263   
  
inv01  �  B�        %� Č +  
,ix221    
  
inv01  �  B�        $dh "� +  
,ix2497   
  
inv01   #� 8� +  
,ix2946   
  
inv01   � �d +  
,ix2978   
  
inv01   �  #� +  
,ix3004   
  
inv01  �  B�        5h s4 +  
,ix2310   
  
inv01   K� �d +  
,ix2340   
  
inv01  �  B�        (k� 8� +  
,ix291    
  
inv01   #�  �� +  
,ix843    
  
inv01  �  B�        ��  +  
,ix2278   
  
inv01   #G@ � +  
,ix913    
  
inv01   $݀ v� +  
,ix1805   
  
inv01  �  B�        &�( � +  
,ix2333   
  
aoi32   *@ �� +  
,ix2782   
  
aoi32   ,�� �T +  
,ix2488   
  
aoi32  �  B�        "�� 
ɸ +  
,ix1856   
  
aoi32  �  B�        �h �� +  
,ix2136   
  
aoi32  �  B�        ,�� �� +  
,ix1704   
  
aoi32  �  B�        $�� Č +  
,ix2638   
  
aoi32  �  B�        % � �� +  
,ix2928   
  
aoi32  �  B�        &9( v� +  
,ix2258   
  
nand02 �  B�        $%� l� +  
,ix3150   
  
nand02  �� l� +  
,ix2072   
  
nand02 �  B�        �( 
ɸ +  
,ix3755   
  
nand02 �  B�        Ҩ tX +  
,ix3324   
  
nand02 �  B�        �( tX +  
,ix3336   
  
nand02  	'� �T +  
,ix3078   
  
nand02  �  �d +  
,ix3068   
  
nand02 �  B�        P� /  +  
,ix2118   
  
nand02  Q� /  +  
,ix2004   
  
nand02 �  B�        h ! +  
,ix2124   
  
nand02 �  B�        *~� /  +  
,ix2824   
  
nand02 �  B�        wh ! +  
,ix2770   
  
nand02  -�  
ɸ +  
,ix2832   
  
nand02  -�  Č +  
,ix2532   
  
nand02  ހ ! +  
,ix2476   
  
nand02 �  B�        �� /  +  
,ix2086   
  
nand02 �  B�        &9( l� +  
,ix1830   
  
nand02 �  B�        �h /  +  
,ix2112   
  
nand02 �  B�        C� %$ +  
,ix1950   
  
nand02  )�  v� +  
,ix2540   
  
nand02  ,O� 
ɸ +  
,ix1748   
  
nand02  Q� �T +  
,ix1692   
  
nand02 �  B�        *@h Č +  
,ix2612   
  
nand02 �  B�        )�� "� +  
,ix1820   
  
nand02  
!� %$ +  
,ix2724   
  
nand02 �  B�        $�( 
ɸ +  
,ix2904   
  
nand02 �  B�        %�� �� +  
,ix2602   
  
nand02 �  B�        "1� /  +  
,ix2082   
  
nand02  Q� #� +  
,ix3016   
  
nand02 �  B�        )� tX +  
,ix2894   
  
nand02  $� /  +  
,ix2104   
  
nand02  *{  l� +  
,ix1756   
  
nand02  �� s4 +  
,ix2352   
  
mux21  �  B�        �< "� +  
,ix3250   
  
mux21   ��  X +  
,ix3399   
  
mux21  �  B�        � l� +  
,ix3353   
  
mux21   !� tX +  
,ix3248   
  
mux21   "�@ l� +  
,ix3371   
  
mux21   !� l� +  
,ix1535   
  
mux21  �  B�        "C| � +  
,ix3134   
  
mux21   �@  X +  
,ix3711   
  
mux21   �   X +  
,ix3468   
  
mux21  �  B�        < "� +  
,ix3382   
  
mux21  �  B�        � "� +  
,ix3641   
  
mux21  �  B�        s|  X +  
,ix3270   
  
mux21   �  "� +  
,ix3361   
  
mux21  �  B�        "�  X +  
,ix3119   
  
mux21   w@  X +  
,ix2056   
  
mux21   %� "� +  
,ix3436   
  
mux21  �  B�        3� "� +  
,ix3703   
  
mux21   �� l� +  
,ix3408   
  
mux21  �  B�        .� l� +  
,ix3379   
  
mux21   �� tX +  
,ix3253   
  
mux21   �  l� +  
,ix3289   
  
mux21   �� "� +  
,ix3727   
  
mux21  �  B�        C< l� +  
,ix3540   
  
mux21   �  � +  
,ix3544   
  
mux21  �  B�        �� tX +  
,ix3735   
  
mux21  �  B�        n| l� +  
,ix3228   
  
mux21   �� tX +  
,ix3447   
  
mux21  �  B�        n| tX +  
,ix3056   
  
mux21  �  B�        
� 
ɸ +  
,ix3463   
  
mux21   <@ � +  
,ix3245   
  
mux21  �  B�        o� 
ɸ +  
,ix3226   
  
mux21  �  B�        �| 
ɸ +  
,ix3209   
  
mux21  �  B�        p� /  +  
,ix1583   
  
mux21  �  B�        �| /  +  
,ix3086   
  
mux21  �  B�        � /  +  
,ix1599   
  
mux21   ;  /  +  
,ix3082   
  
mux21  �  B�        �� � +  
,ix3217   
  
mux21  �  B�        �< tX +  
,ix3167   
  
mux21  �  B�        �� tX +  
,ix2008   
  
mux21   �� � +  
,ix3183   
  
mux21   l@ � +  
,ix1958   
  
mux21  �  B�        I< tX +  
,ix3294   
  
mux21  �  B�        �|  X +  
,ix3328   
  
mux21   �@ "� +  
,ix3529   
  
mux21   �  X +  
,ix3358   
  
mux21   �� "� +  
,ix3585   
  
mux21  �  B�        E�  X +  
,ix3242   
  
mux21  �  B�        2| "� +  
,ix3415   
  
mux21  �  B�        � l� +  
,ix3234   
  
mux21  �  B�        	� l� +  
,ix3431   
  
mux21  �  B�        
�  X +  
,ix3719   
  
mux21   
�  "� +  
,ix3500   
  
mux21   J� tX +  
,ix3317   
  
mux21   @ � +  
,ix3240   
  
mux21   ̀ � +  
,ix3281   
  
mux21  �  B�         n� � +  
,ix1551   
  
mux21  �  B�        a| 
ɸ +  
,ix3118   
  
mux21  �  B�        �� 
ɸ +  
,ix1567   
  
mux21   �� 
ɸ +  
,ix3102   
  
mux21  �  B�        X� "� +  
,ix3278   
  
mux21   @  X +  
,ix3325   
  
mux21  �  B�        ��  X +  
,ix3135   
  
mux21  �  B�        |  X +  
,ix2040   
  
mux21  �  B�        ~< l� +  
,ix3151   
  
mux21  �  B�        �< l� +  
,ix2024   
  
mux21   �� l� +  
,ix3286   
  
mux21  �  B�        ڼ 
ɸ +  
,ix3232   
  
mux21   )�  tX +  
,ix1231   
  
mux21   ,�� tX +  
,ix1133   
  
mux21  �  B�        '%| l� +  
,ix3158   
  
mux21   !r� �� +  
,ix2874   
  
mux21  �  B�         O| Č +  
,ix3044   
  
mux21   @  v� +  
,ix1431   
  
mux21  �  B�        (�| � +  
,ix3050   
  
mux21   -i  � +  
,ix2880   
  
mux21   '�  tX +  
,ix1483   
  
mux21   %�@ 
ɸ +  
,ix1239   
  
mux21  �  B�        )W� 
ɸ +  
,ix1141   
  
mux21   $݀ 
ɸ +  
,ix3174   
  
mux21  �  B�        �| �T +  
,ix1247   
  
mux21   �� Č +  
,ix1149   
  
mux21   �  Č +  
,ix3190   
  
mux21   C� �T +  
,ix2866   
  
mux21  �  B�        ¼ �T +  
,ix3038   
  
mux21   h� Č +  
,ix1379   
  
mux21  �  B�        P| �T +  
,ix3072   
  
mux21  �  B�        	��  +  
,ix1263   
  
mux21  �  B�        	�� 8� +  
,ix1165   
  
mux21  �  B�        ]�  +  
,ix1255   
  
mux21   a�  +  
,ix1157   
  
mux21     Č +  
,ix3206   
  
mux21   T@ 8� +  
,ix2856   
  
mux21   y� 8� +  
,ix3032   
  
mux21   T@ �T +  
,ix1327   
  
mux21   C� #� +  
,ix2564   
  
mux21  �  B�         | %$ +  
,ix2740   
  
mux21  �  B�        9� #� +  
,ix1315   
  
mux21  �  B�        | ! +  
,ix3060   
  
mux21     #� +  
,ix641    
  
mux21  �  B�        ?� ! +  
,ix543    
  
mux21   @ %$ +  
,ix633    
  
mux21  �  B�        �� %$ +  
,ix535    
  
mux21   �@ #� +  
,ix3096   
  
mux21  �  B�         �< #� +  
,ix2574   
  
mux21   "M@ %$ +  
,ix2746   
  
mux21   � #� +  
,ix1367   
  
mux21   #�  #� +  
,ix625    
  
mux21   %y� #� +  
,ix527    
  
mux21   #�� ! +  
,ix3112   
  
mux21   (�@ ! +  
,ix2580   
  
mux21  �  B�        &+| ! +  
,ix2752   
  
mux21   "�  ! +  
,ix1419   
  
mux21  �  B�        �< �� +  
,ix2225   
  
mux21   �  �� +  
,ix2127   
  
mux21  �  B�        � Č +  
,ix2217   
  
mux21  �  B�        � Č +  
,ix2119   
  
mux21   m� v� +  
,ix2416   
  
mux21   l@ /  +  
,ix2438   
  
mux21   �� Č +  
,ix2202   
  
mux21  �  B�        �� �T +  
,ix2444   
  
mux21  �  B�        
7< Č +  
,ix2911   
  
mux21   �@ �� +  
,ix2212   
  
mux21  �  B�        >| Č +  
,ix2422   
  
mux21   �@ /  +  
,ix2963   
  
mux21   |  v� +  
,ix2209   
  
mux21  �  B�        r< �� +  
,ix2111   
  
mux21  �  B�        �< /  +  
,ix2394   
  
mux21  �  B�        !� v� +  
,ix2220   
  
mux21  �  B�        @� /  +  
,ix2400   
  
mux21   �� � +  
,ix3015   
  
mux21   R  l� +  
,ix2092   
  
mux21   F  tX +  
,ix2193   
  
mux21  �  B�        �� tX +  
,ix2095   
  
mux21  �  B�        �� 
ɸ +  
,ix2201   
  
mux21   �� � +  
,ix2103   
  
mux21  �  B�        �| tX +  
,ix2374   
  
mux21   R  � +  
,ix2380   
  
mux21  �  B�        H< � +  
,ix2228   
  
mux21  �  B�        �< tX +  
,ix3067   
  
mux21   '��  X +  
,ix2717   
  
mux21   #�   X +  
,ix2066   
  
mux21   �  � +  
,ix1798   
  
mux21   �@ 
ɸ +  
,ix1982   
  
mux21   �  l� +  
,ix3003   
  
mux21  �  B�        z� "� +  
,ix2823   
  
mux21   �� "� +  
,ix2725   
  
mux21   ,�  X +  
,ix2050   
  
mux21  �  B�        !*< "� +  
,ix1988   
  
mux21   !�@  X +  
,ix1806   
  
mux21   ��  X +  
,ix3055   
  
mux21  �  B�        �� v� +  
,ix2831   
  
mux21   �@ v� +  
,ix2733   
  
mux21   I� /  +  
,ix2034   
  
mux21   �  v� +  
,ix2839   
  
mux21   	�� �� +  
,ix2741   
  
mux21   
�� v� +  
,ix2018   
  
mux21     �� +  
,ix1790   
  
mux21   B@ v� +  
,ix1976   
  
mux21   t� /  +  
,ix2951   
  
mux21  �  B�        t| �� +  
,ix1780   
  
mux21   E� Č +  
,ix1970   
  
mux21  �  B�        �< v� +  
,ix2899   
  
mux21  �  B�        �| v� +  
,ix1996   
  
mux21  �  B�        "� �� +  
,ix2749   
  
mux21  �  B�        "� v� +  
,ix2847   
  
mux21   '   X +  
,ix2815   
  
mux21  �  B�        o� s4 +  
,ix2162   
  
mux21  �  B�        �� �T +  
,ix2168   
  
mux21   @ �T +  
,ix1751   
  
mux21   �  s4 +  
,ix1759   
  
mux21   e@ /  +  
,ix1735   
  
mux21   ,O� 8� +  
,ix693    
  
mux21  �  B�        � s4 +  
,ix701    
  
mux21   �� ! +  
,ix805    
  
mux21  �  B�         0< �d +  ,ix79   
  
mux21   %� v� +  
,ix1743   
  
mux21  �  B�        %P� s4 +  
,ix2778   
  
mux21  �  B�        -?� �d +  
,ix2484   
  
mux21   p  �d +  
,ix2774   
  
mux21  �  B�        �� ! +  
,ix2480   
  
mux21   $@ s4 +  
,ix2808   
  
mux21   &T� s4 +  
,ix2814   
  
mux21  �  B�        a| s4 +  
,ix789    
  
mux21  �  B�        �| s4 +  
,ix797    
  
mux21   -I� �d +  ,ix71   
  
mux21   �@ ! +  
,ix183    
  
mux21  �  B�        "� 8� +  
,ix2389   
  
mux21  �  B�        - � /  +  
,ix773    
  
mux21   *{  8� +  
,ix781    
  
mux21  �  B�        ��  +  
,ix2285   
  
mux21   "�   +  
,ix1700   
  
mux21   0@  +  
,ix1696   
  
mux21   2� ! +  
,ix243    
  
mux21  �  B�        /� %$ +  
,ix2553   
  
mux21   � 8� +  
,ix2449   
  
mux21   !�� v� +  
,ix2441   
  
mux21   �  �� +  
,ix1655   
  
mux21   >� �d +  
,ix1663   
  
mux21  �  B�        �| #� +  
,ix1767   
  
mux21  �  B�        H< 8� +  
,ix1892   
  
mux21  �  B�        "�� s4 +  
,ix2670   
  
mux21   ��  +  
,ix2132   
  
mux21  �  B�        �| �d +  
,ix1924   
  
mux21  �  B�        �� %$ +  
,ix2700   
  
mux21  �  B�        	�� ! +  
,ix2128   
  
mux21  �  B�        �� #� +  
,ix2516   
  
mux21   *�  ! +  
,ix2522   
  
mux21    �@ ! +  
,ix167    
  
mux21  �  B�        4� #� +  
,ix175    
  
mux21   �  8� +  
,ix1923   
  
mux21   �@ 8� +  
,ix2320   
  
mux21  �  B�        R� 8� +  
,ix1915   
  
mux21   �� �T +  
,ix2288   
  
mux21   �� �� +  
,ix1907   
  
mux21  �  B�        !�< /  +  
,ix1899   
  
mux21  �  B�        &Ǽ  +  
,ix2277   
  
mux21   +U� Č +  
,ix151    
  
mux21   *�  s4 +  
,ix159    
  
mux21   �� �d +  
,ix865    
  
mux21  �  B�        %1| 8� +  
,ix857    
  
mux21  �  B�        �� %$ +  
,ix347    
  
mux21  �  B�        "�� �T +  
,ix235    
  
mux21  �  B�        � #� +  
,ix2545   
  
mux21  �  B�        �< �d +  
,ix1918   
  
mux21   P� 8� +  
,ix2537   
  
mux21   ��  +  
,ix1886   
  
mux21    � tX +  
,ix2529   
  
mux21  �  B�        ( < "� +  
,ix2521   
  
mux21    �@ s4 +  
,ix2962   
  
mux21  �  B�        �< #� +  
,ix2992   
  
mux21  �  B�        (>� �� +  
,ix609    
  
mux21  �  B�        *| �� +  
,ix511    
  
mux21   %�  /  +  
,ix3144   
  
mux21  �  B�        (�| �d +  
,ix617    
  
mux21   )�@ �d +  
,ix519    
  
mux21   )#@ s4 +  
,ix3128   
  
mux21  �  B�        )�|  +  
,ix2758   
  
mux21  �  B�        *�< �T +  
,ix2588   
  
mux21   'N� �T +  
,ix1471   
  
mux21  �  B�        5� #� +  
,ix969    
  
mux21   � %$ +  
,ix339    
  
mux21  �  B�        [| %$ +  
,ix2694   
  
mux21   � ! +  
,ix331    
  
mux21  �  B�        #�� �d +  
,ix2664   
  
mux21   %�� �d +  
,ix323    
  
mux21  �  B�        ( < Č +  
,ix315    
  
mux21  �  B�        �� �d +  
,ix1931   
  
mux21   �  s4 +  
,ix1827   
  
mux21   �@ �T +  
,ix1819   
  
mux21   F  8� +  
,ix2294   
  
mux21   �@ �d +  
,ix2326   
  
mux21  �  B�        �� ! +  
,ix961    
  
mux21  �  B�        �� 8� +  
,ix2986   
  
mux21  �  B�        � 8� +  
,ix953    
  
mux21    �@  +  
,ix2956   
  
mux21  �  B�        %P� �T +  
,ix945    
  
mux21  �  B�        )w< � +  
,ix937    
  
mux21  �  B�        j� �T +  
,ix1732   
  
mux21   @ Č +  
,ix1738   
  
mux21  �  B�        | Č +  
,ix2373   
  
mux21  �  B�        �<  +  
,ix2381   
  
mux21  �  B�        +�� tX +  
,ix2357   
  
mux21  �  B�        #�< �� +  
,ix2365   
  nor02ii  �  B�        B� l� +  
,ix3383   
  nor02ii   �� v� +  
,ix3909   
  nor02ii  �  B�        �� �� +  
,ix3911   
  nor02ii  �  B�        �� 
ɸ +  
,ix3479   
  nor02ii  �  B�        ,r� l� +  
,ix2888   
  nor02ii   +@ l� +  
,ix3054   
  nor02ii  �  B�        
d( �T +  
,ix1269   
  nor02ii   �� 8� +  
,ix647    
  nor02ii  �  B�        �� /  +  
,ix2231   
  nor02ii   �@ � +  
,ix2078   
  nor02ii   &� � +  
,ix2088   
  nor02ii   -�  #� +  ,ix9    
  nor02ii   *{   X +  
,ix1814   
  nor02ii   )��  X +  
,ix1992   
  nor02ii  �  B�        �� 
ɸ +  
,ix2853   
  nor02ii   � s4 +  
,ix1777   
  nor02ii   Y  s4 +  
,ix2356   
  nor02ii   /  �d +  
,ix815    
  nor02ii   y� �d +  
,ix3020   
  nor02ii   6@ ! +  
,ix193    
  nor02ii   z� ! +  
,ix2728   
  nor02ii   @ %$ +  
,ix2563   
  nor02ii  �  B�        �� %$ +  
,ix1946   
  nor02ii   K�  +  
,ix2399   
  nor02ii  �  B�        �( �T +  
,ix1954   
  nor02ii   H@ %$ +  
,ix357    
  nor02ii  �  B�        ,� %$ +  
,ix2720   
  nor02ii  �  B�        (�( v� +  
,ix2596   
  nor02ii  �  B�        '� v� +  
,ix2762   
  nor02ii   @ ! +  
,ix979    
  nor02ii  �  B�        �� ! +  
,ix3012   
  nor02ii  �  B�        �� 8� +  
,ix1941   
  nor02ii    � �T +  
,ix2348   
  
oai21   *�@ /  +  
,ix2830   
  
oai21   ,�@ l� +  
,ix2890   
  
oai21  �  B�        -ʨ Č +  
,ix2538   
  
oai21  �  B�        �h 
ɸ +  
,ix2084   
  
oai21  �  B�        &� "� +  
,ix1828   
  
oai21   �� /  +  
,ix2110   
  
oai21  �  B�        )e� v� +  
,ix2598   
  
oai21  �  B�        ,4h 
ɸ +  
,ix1754   
  
oai21  �  B�        (�( Č +  
,ix2610   
  
oai21   )�@ "� +  
,ix1818   
  
oai21   %�  � +  
,ix2902   
  
oai21   %�@ �� +  
,ix2600   
  
oai21  �  B�         �� 
ɸ +  
,ix2080   
  
oai21   )�� l� +  
,ix2892   
  
oai21  �  B�        #�h /  +  
,ix2102   
  
oai21   *[� "� +  
,ix1816   
  
aoi22   >� /  +  
,ix2174   
  
aoi22  �  B�        ,Ш v� +  
,ix2820   
  
aoi22  �  B�        ,S�  +  
,ix2528   
  
aoi22  �  B�        $� v� +  
,ix2250   
  
aoi22  �  B�        #�h "� +  
,ix1848   
  
aoi22   '/@ 8� +  
,ix2630   
  
aoi22   $�@ � +  
,ix2920   
  
aoi22  �  B�        &w� tX +  
,ix1744   
  
xnor2  �  B�        X #� +  
,ix3590   
  
xnor2   #  Č +  
,ix3799   
  
xnor2  �  B�        u� �� +  
,ix3795   
  
xnor2   ��  X +  
,ix3791   
  
xnor2  �  B�        �X  X +  
,ix3787   
  
xnor2  �  B�        G�  X +  
,ix3783   
  
xnor2  �  B�        G� "� +  
,ix3779   
  
xnor2  �  B�        A� l� +  
,ix3775   
  
xnor2   � /  +  
,ix3767   
  
xnor2  �  B�        � /  +  
,ix3759   
  
xnor2   �  "� +  
,ix3264   
  
xnor2  �  B�        !� l� +  
,ix3156   
  
xnor2   #�@ tX +  
,ix3164   
  
xnor2  �  B�        � "� +  
,ix3596   
  
xnor2   O�  X +  
,ix3272   
  
xnor2   �   X +  
,ix3466   
  
xnor2  �  B�        �X l� +  
,ix3578   
  
xnor2   ��  X +  
,ix3268   
  
xnor2   �  "� +  
,ix3643   
  
xnor2   }@  X +  
,ix2362   
  
xnor2   �� "� +  
,ix2090   
  
xnor2   �� "� +  
,ix3434   
  
xnor2   �� "� +  
,ix3801   
  
xnor2   �� l� +  
,ix3588   
  
xnor2   �  l� +  
,ix2392   
  
xnor2  �  B�        � � +  
,ix3614   
  
xnor2  �  B�        �� 
ɸ +  
,ix3300   
  
xnor2  �  B�        G� 
ɸ +  
,ix3320   
  
xnor2  �  B�        G� l� +  
,ix3554   
  
xnor2  �  B�        �� "� +  
,ix3608   
  
xnor2  �  B�        nX l� +  
,ix3288   
  
xnor2   x@ "� +  
,ix3538   
  
xnor2  �  B�        �� � +  
,ix3296   
  
xnor2  �  B�        �� tX +  
,ix3292   
  
xnor2   z� /  +  
,ix3204   
  
xnor2   s� v� +  
,ix3212   
  
xnor2   y� v� +  
,ix3220   
  
xnor2  �  B�        �� � +  
,ix2436   
  
xnor2  �  B�        
� 
ɸ +  
,ix2448   
  
xnor2   �� tX +  
,ix2426   
  
xnor2  �  B�        
� /  +  
,ix3222   
  
xnor2   �  tX +  
,ix2414   
  
xnor2  �  B�        �  X +  
,ix3562   
  
xnor2  �  B�        
� l� +  
,ix3284   
  
xnor2   �@ "� +  
,ix3531   
  
xnor2   ��  X +  
,ix3570   
  
xnor2   <@ "� +  
,ix3276   
  
xnor2  �  B�        � "� +  
,ix3587   
  
xnor2   
!�  X +  
,ix3602   
  
xnor2   �� l� +  
,ix3280   
  
xnor2   	�  "� +  
,ix3498   
  
xnor2    x� � +  
,ix3172   
  
xnor2  �  B�        aX 
ɸ +  
,ix3180   
  
xnor2   �� 
ɸ +  
,ix3188   
  
xnor2   $@  X +  
,ix2382   
  
xnor2   ��  X +  
,ix2372   
  
xnor2   �  l� +  
,ix2404   
  
xnor2   ƀ 
ɸ +  
,ix3196   
  
xnor2  �  B�         t� �� +  
,ix3186   
  
xnor2    x� �� +  
,ix3184   
  
xnor2  �  B�        -e � +  
,ix1095   
  
xnor2  �  B�        )]� tX +  
,ix3170   
  
xnor2   -�@ tX +  
,ix3168   
  
xnor2  �  B�        (� 
ɸ +  
,ix1083   
  
xnor2   &�  
ɸ +  
,ix1447   
  
xnor2   )a� 
ɸ +  
,ix1453   
  
xnor2   �@ �T +  
,ix1059   
  
xnor2  �  B�        �� Č +  
,ix1395   
  
xnor2   �� Č +  
,ix1401   
  
xnor2  �  B�         �T +  
,ix1047   
  
xnor2  �  B�        d� Č +  
,ix3202   
  
xnor2   C� Č +  
,ix3200   
  
xnor2  �  B�        
��  +  
,ix1291   
  
xnor2   
� 8� +  
,ix1297   
  
xnor2  �  B�        �� 8� +  
,ix1003   
  
xnor2  �  B�        ]�  +  
,ix1035   
  
xnor2  �  B�        � �T +  
,ix1343   
  
xnor2  �  B�        � �T +  
,ix1349   
  
xnor2  �  B�        o� s4 +  
,ix1023   
  
xnor2  �  B�        ��  +  
,ix3218   
  
xnor2   ��  +  
,ix3216   
  
xnor2  �  B�        ,�� tX +  
,ix1107   
  
xnor2   ()@ l� +  
,ix1499   
  
xnor2  �  B�        (%X l� +  
,ix1505   
  
xnor2  �  B�        !�X Č +  
,ix1071   
  
xnor2  �  B�        %V� ! +  
,ix3124   
  
xnor2   '�@ ! +  
,ix3122   
  
xnor2  �  B�        K� %$ +  
,ix401    
  
xnor2  �  B�         X %$ +  
,ix3092   
  
xnor2   $@ %$ +  
,ix3090   
  
xnor2  �  B�        d� #� +  
,ix1279   
  
xnor2   $@ ! +  
,ix1285   
  
xnor2  �  B�         #� +  
,ix381    
  
xnor2  �  B�        � %$ +  
,ix413    
  
xnor2  �  B�        � %$ +  
,ix1331   
  
xnor2   �� %$ +  
,ix1337   
  
xnor2    �@ %$ +  
,ix425    
  
xnor2   !�  #� +  
,ix3108   
  
xnor2    �  #� +  
,ix3106   
  
xnor2  �  B�        #� #� +  
,ix437    
  
xnor2   $� #� +  
,ix1383   
  
xnor2   &T� #� +  
,ix1389   
  
xnor2  �  B�        '�X ! +  
,ix449    
  
xnor2  �  B�        �� Č +  
,ix2875   
  
xnor2   �� �� +  
,ix2881   
  
xnor2   S   +  
,ix1985   
  
xnor2   -� �T +  
,ix2432   
  
xnor2   l@ Č +  
,ix2430   
  
xnor2   �  �T +  
,ix2009   
  
xnor2  �  B�        >X v� +  
,ix2410   
  
xnor2   �  �� +  
,ix2408   
  
xnor2   |  �� +  
,ix2021   
  
xnor2   V� v� +  
,ix2979   
  
xnor2  �  B�        x v� +  
,ix2985   
  
xnor2   �  �� +  
,ix2033   
  
xnor2  �  B�        � 
ɸ +  
,ix2388   
  
xnor2  �  B�        �� � +  
,ix2386   
  
xnor2   &� l� +  
,ix3083   
  
xnor2   ,� l� +  
,ix3089   
  
xnor2    � tX +  
,ix2069   
  
xnor2   �� 
ɸ +  
,ix2045   
  
xnor2  �  B�        �� � +  
,ix3031   
  
xnor2   �� � +  
,ix3037   
  
xnor2   ,� � +  
,ix2057   
  
xnor2   �  tX +  
,ix2368   
  
xnor2  �  B�        � tX +  
,ix2366   
  
xnor2  �  B�        � Č +  
,ix1965   
  
xnor2  �  B�        7 Č +  
,ix1997   
  
xnor2  �  B�        JX �� +  
,ix2927   
  
xnor2  �  B�        DX �� +  
,ix2933   
  
xnor2  �  B�        ��  X +  
,ix3019   
  
xnor2   �  X +  
,ix3025   
  
xnor2  �  B�        "* "� +  
,ix2679   
  
xnor2    �@  X +  
,ix2062   
  
xnor2   "�   X +  
,ix2060   
  
xnor2  �  B�        �X �� +  
,ix2643   
  
xnor2  �  B�        E� /  +  
,ix2967   
  
xnor2   $@ /  +  
,ix2973   
  
xnor2   �� �� +  
,ix2619   
  
xnor2  �  B�        	�� v� +  
,ix2915   
  
xnor2   	�� v� +  
,ix2921   
  
xnor2  �  B�         �� +  
,ix2631   
  
xnor2  �  B�         v� +  
,ix2030   
  
xnor2  �  B�         v� +  
,ix2028   
  
xnor2   �� �T +  
,ix2607   
  
xnor2   �  v� +  
,ix2014   
  
xnor2  �  B�        �X v� +  
,ix2012   
  
xnor2  �  B�        "� v� +  
,ix2863   
  
xnor2   �� �� +  
,ix2869   
  
xnor2  �  B�        �� Č +  
,ix2587   
  
xnor2   (ŀ  X +  
,ix2691   
  
xnor2  �  B�        %u�  X +  
,ix3071   
  
xnor2  �  B�        &o�  X +  
,ix3077   
  
xnor2   v  /  +  
,ix2655   
  
xnor2  �  B�        R� l� +  
,ix2046   
  
xnor2   V� l� +  
,ix2044   
  
xnor2   _@ "� +  
,ix2667   
  
xnor2  �  B�        + �d +  
,ix2860   
  
xnor2   	�� �d +  
,ix1673   
  
xnor2  �  B�        )� ! +  
,ix2206   
  
xnor2   �  s4 +  
,ix1977   
  
xnor2   �� s4 +  
,ix1015   
  
xnor2  �  B�        ��  +  
,ix2005   
  
xnor2  �  B�        � Č +  
,ix2029   
  
xnor2  �  B�        X �T +  
,ix2017   
  
xnor2   	�� s4 +  
,ix1993   
  
xnor2   e@ 
ɸ +  
,ix2065   
  
xnor2  �  B�        l �d +  
,ix717    
  
xnor2  �  B�        &P� s4 +  
,ix733    
  
xnor2   *�@ v� +  
,ix2838   
  
xnor2   +U� 8� +  
,ix2818   
  
xnor2  �  B�        �� s4 +  
,ix2812   
  
xnor2   � ! +  
,ix2806   
  
xnor2   8� #� +  ,ix95   
  
xnor2   ,�� ! +  
,ix111    
  
xnor2   !4  �d +  
,ix2520   
  
xnor2   �� 
ɸ +  
,ix2230   
  
xnor2    @ v� +  
,ix2041   
  
xnor2   )  /  +  
,ix2826   
  
xnor2  �  B�        aX /  +  
,ix1725   
  
xnor2   -�� 8� +  
,ix2788   
  
xnor2  �  B�        �� /  +  
,ix1713   
  
xnor2  �  B�        ${� s4 +  
,ix2790   
  
xnor2  �  B�        !� v� +  
,ix1705   
  
xnor2  �  B�        @� s4 +  
,ix2794   
  
xnor2  �  B�        ��  +  
,ix2190   
  
xnor2   J� �d +  
,ix2796   
  
xnor2  �  B�        ��  +  
,ix1689   
  
xnor2  �  B�        � ! +  
,ix2800   
  
xnor2   
� �d +  
,ix2196   
  
xnor2  �  B�        ,k �d +  
,ix2498   
  
xnor2   '/@ s4 +  
,ix2844   
  
xnor2   �@ s4 +  
,ix2502   
  
xnor2  �  B�        �� s4 +  
,ix727    
  
xnor2  �  B�        � ! +  
,ix2504   
  
xnor2   �  s4 +  
,ix2850   
  
xnor2  �  B�        X ! +  
,ix2508   
  
xnor2  �  B�        �� s4 +  
,ix711    
  
xnor2  �  B�        ژ ! +  
,ix2568   
  
xnor2  �  B�        �� #� +  
,ix393    
  
xnor2  �  B�         X s4 +  
,ix1043   
  
xnor2   &5@ 8� +  
,ix1067   
  
xnor2   k@ s4 +  
,ix1055   
  
xnor2   �@ s4 +  
,ix1031   
  
xnor2   ,�� s4 +  
,ix2526   
  
xnor2   �  ! +  
,ix2514   
  
xnor2  �  B�        "� 8� +  
,ix1730   
  
xnor2  �  B�        -� 
ɸ +  
,ix1103   
  
xnor2   -I� /  +  
,ix2882   
  
xnor2   *[� Č +  
,ix1079   
  
xnor2   -�� �T +  
,ix2546   
  
xnor2   6@  +  
,ix2301   
  
xnor2  �  B�        "�  +  
,ix2317   
  
xnor2  �  B�        ��  +  
,ix1736   
  
xnor2  �  B�        ,K� /  +  
,ix763    
  
xnor2  �  B�        +� �T +  
,ix2534   
  
xnor2   ,�  v� +  
,ix751    
  
xnor2   -�� s4 +  
,ix2496   
  
xnor2  �  B�        *w 8� +  
,ix743    
  
xnor2  �  B�        �� %$ +  
,ix1926   
  
xnor2  �  B�        	�X #� +  
,ix2154   
  
xnor2  �  B�        �� %$ +  
,ix1934   
  
xnor2  �  B�        � #� +  
,ix2605   
  
xnor2   � ! +  
,ix2668   
  
xnor2   �� %$ +  
,ix1922   
  
xnor2   %� 8� +  
,ix1890   
  
xnor2    �@ 
ɸ +  
,ix1854   
  
xnor2   �� %$ +  
,ix259    
  
xnor2  �  B�        #�� s4 +  
,ix275    
  
xnor2   
� ! +  
,ix1679   
  
xnor2  �  B�        ��  +  
,ix1695   
  
xnor2  �  B�        � /  +  
,ix2184   
  
xnor2   �  �� +  
,ix2172   
  
xnor2  �  B�        :� �d +  
,ix2166   
  
xnor2  �  B�        	#� ! +  
,ix2160   
  
xnor2  �  B�        �X �d +  
,ix2465   
  
xnor2   R  8� +  
,ix2481   
  
xnor2   $�@ l� +  
,ix1840   
  
xnor2   #G@ 
ɸ +  
,ix1842   
  
xnor2  �  B�        gX v� +  
,ix2178   
  
xnor2  �  B�        "�X Č +  
,ix1862   
  
xnor2  �  B�        � �� +  
,ix2142   
  
xnor2   L  8� +  
,ix1878   
  
xnor2   k@  +  
,ix2144   
  
xnor2  �  B�        !� 8� +  
,ix1894   
  
xnor2   � �d +  
,ix2148   
  
xnor2  �  B�        �� �d +  
,ix1910   
  
xnor2  �  B�        	�� �d +  
,ix2150   
  
xnor2  �  B�         8� +  
,ix1718   
  
xnor2    :  �d +  
,ix105    
  
xnor2   \� 8� +  
,ix1853   
  
xnor2      +  
,ix1720   
  
xnor2  �  B�        (� #� +  
,ix2558   
  
xnor2  �  B�        &X s4 +  
,ix2304   
  
xnor2  �  B�        �� s4 +  
,ix1724   
  
xnor2  �  B�        ` #� +  ,ix89   
  
xnor2  �  B�        U s4 +  
,ix1837   
  
xnor2   Q�  +  
,ix1784   
  
xnor2   @  +  
,ix2599   
  
xnor2  �  B�        �� #� +  
,ix421    
  
xnor2  �  B�        *� ! +  
,ix445    
  
xnor2   !�  ! +  
,ix433    
  
xnor2   >� #� +  
,ix409    
  
xnor2   �� 8� +  
,ix1995   
  
xnor2  �  B�        �X 8� +  
,ix2007   
  
xnor2  �  B�        X �T +  
,ix2019   
  
xnor2   �  Č +  
,ix2031   
  
xnor2  �  B�        �� �� +  
,ix2043   
  
xnor2  �  B�         �X /  +  
,ix2067   
  
xnor2  �  B�        'J� �T +  
,ix1742   
  
xnor2   +@ �� +  
,ix481    
  
xnor2   *�@  +  
,ix2590   
  
xnor2  �  B�        +q �d +  
,ix457    
  
xnor2  �  B�        aX v� +  
,ix2236   
  
xnor2  �  B�        +Q� 
ɸ +  
,ix1762   
  
xnor2   ,0� Č +  
,ix141    
  
xnor2   "M@ /  +  
,ix1889   
  
xnor2   -�@ �� +  
,ix1750   
  
xnor2   ,o   +  
,ix129    
  
xnor2    �� v� +  
,ix1877   
  
xnor2  �  B�        'ǘ  +  
,ix1712   
  
xnor2   +�� s4 +  
,ix121    
  
xnor2   �� �� +  
,ix1869   
  
xnor2   #��  +  
,ix1714   
  
xnor2   +�� ! +  
,ix2552   
  
xnor2   �� �T +  
,ix2272   
  
xnor2    �� tX +  
,ix2491   
  
xnor2   8� ! +  
,ix2672   
  
xnor2   q@  +  
,ix1870   
  
xnor2  �  B�        �� %$ +  
,ix2686   
  
xnor2  �  B�        F� s4 +  
,ix2475   
  
xnor2   
�@ #� +  
,ix2702   
  
xnor2   �  �d +  
,ix1902   
  
xnor2  �  B�        
� %$ +  
,ix2710   
  
xnor2  �  B�        /� #� +  
,ix2459   
  
xnor2   ހ %$ +  
,ix399    
  
xnor2   e@ �d +  
,ix2960   
  
xnor2  �  B�        %u�  +  
,ix2926   
  
xnor2  �  B�        �� %$ +  
,ix2698   
  
xnor2   #�� �T +  
,ix2636   
  
xnor2  �  B�        �� �d +  
,ix2617   
  
xnor2  �  B�        ,X s4 +  
,ix2629   
  
xnor2   ��  +  
,ix2641   
  
xnor2  �  B�        �X v� +  
,ix2653   
  
xnor2   �� l� +  
,ix2665   
  
xnor2   (
  "� +  
,ix2689   
  
xnor2   �  #� +  
,ix881    
  
xnor2    �� 8� +  
,ix897    
  
xnor2   (ŀ Č +  
,ix2622   
  
xnor2  �  B�        #$ "� +  
,ix1834   
  
xnor2   %;@ Č +  
,ix2624   
  
xnor2  �  B�        '+X "� +  
,ix2511   
  
xnor2   "�� �T +  
,ix2642   
  
xnor2   $� "� +  
,ix2499   
  
xnor2   "� 8� +  
,ix2656   
  
xnor2   �� ! +  
,ix1021   
  
xnor2  �  B�        5� #� +  
,ix2990   
  
xnor2   @ %$ +  
,ix411    
  
xnor2   _@ %$ +  
,ix423    
  
xnor2   �@ ! +  
,ix435    
  
xnor2  �  B�        $�� �d +  
,ix447    
  
xnor2   &р �d +  
,ix459    
  
xnor2  �  B�        'i� �� +  
,ix483    
  
xnor2  �  B�        �� �d +  
,ix2324   
  
xnor2   V� 8� +  
,ix2292   
  
xnor2   �� Č +  
,ix2256   
  
xnor2   #�@ � +  
,ix2914   
  
xnor2   'ˀ  +  
,ix2616   
  
xnor2  �  B�        �X �d +  
,ix1843   
  
xnor2  �  B�        �X �T +  
,ix1859   
  
xnor2  �  B�        $٘ v� +  
,ix2916   
  
xnor2  �  B�        '+X Č +  
,ix305    
  
xnor2   %;@ 8� +  
,ix2934   
  
xnor2   (�  8� +  
,ix293    
  
xnor2   !� 8� +  
,ix2948   
  
xnor2  �  B�        %�� �d +  
,ix285    
  
xnor2  �  B�        	� �d +  
,ix2964   
  
xnor2  �  B�        #$ �d +  
,ix2650   
  
xnor2  �  B�        �X #� +  
,ix2980   
  
xnor2  �  B�        �� ! +  
,ix269    
  
xnor2   	�@ #� +  
,ix2994   
  
xnor2   e@ %$ +  
,ix2680   
  
xnor2   Q� ! +  
,ix3000   
  
xnor2  �  B�        �� %$ +  
,ix253    
  
xnor2  �  B�        )>� �� +  
,ix485    
  
xnor2  �  B�        'i� /  +  
,ix1487   
  
xnor2   (
  /  +  
,ix1493   
  
xnor2  �  B�        )�X �d +  
,ix461    
  
xnor2  �  B�        )X s4 +  
,ix1435   
  
xnor2   )�  s4 +  
,ix1441   
  
xnor2   )�@  +  
,ix473    
  
xnor2  �  B�        )X �T +  
,ix3140   
  
xnor2  �  B�        *X �T +  
,ix3138   
  
xnor2   �  Č +  
,ix1768   
  
xnor2   e@ s4 +  
,ix891    
  
xnor2   |  �d +  
,ix2312   
  
xnor2   @ �T +  
,ix2311   
  
xnor2  �  B�        % 8� +  
,ix2972   
  
xnor2  �  B�        G� �d +  
,ix2328   
  
xnor2  �  B�        2X  +  
,ix1774   
  
xnor2   �� �d +  
,ix875    
  
xnor2  �  B�        �� s4 +  
,ix2336   
  
xnor2   @  +  
,ix2295   
  
xnor2  �  B�        � 8� +  
,ix1983   
  
xnor2  �  B�        �� �d +  
,ix1033   
  
xnor2  �  B�        �� 8� +  
,ix1045   
  
xnor2   �� 8� +  
,ix1057   
  
xnor2    �  �T +  
,ix1069   
  
xnor2  �  B�        %� /  +  
,ix1081   
  
xnor2  �  B�        *w � +  
,ix1105   
  
xnor2  �  B�        �� Č +  
,ix2627   
  
xnor2  �  B�        l �� +  
,ix2651   
  
xnor2   @ Č +  
,ix2639   
  
xnor2  �  B�        � �T +  
,ix2615   
  
xnor2   &р � +  
,ix2908   
  
xnor2  �  B�        #ߘ v� +  
,ix2242   
  
xnor2  �  B�        ,X "� +  
,ix2687   
  
xnor2  �  B�        %�X tX +  
,ix1808   
  
xnor2  �  B�        #�X tX +  
,ix2663   
  
xnor2   *{  � +  
,ix927    
  
xnor2   &T� v� +  
,ix2244   
  
xnor2   +u  � +  
,ix2347   
  
xnor2  �  B�        #CX � +  
,ix915    
  
xnor2  �  B�        [X  +  
,ix2264   
  
xnor2   &�  tX +  
,ix2335   
  
xnor2   %Z� �T +  
,ix907    
  
xnor2   �  �T +  
,ix2280   
  
xnor2  �  B�        #�X Č +  
,ix2327   
  
xnor2  �  B�         �X  +  
,ix2942   
  
xnor2  �  B�        ��  +  
,ix2296   
  via4  | T   
  via3  |    
  via3   
ϔ   
  via2  � ��   
  via3  �$ ��   
  via3  �$ #CX   
  via2  bx #۰   
  via3  *B\ �l   
  via2  *X 	��   
  via3  )�H 	��   
  via2  (�0 ��   
  via3  )�  �h   
  via2  )�H ��   
  via3  &� �T   
  via3  %�� sX   
  via3  &� �,   
  via2  �X 6�   
  via3  ?, 6�   
  via3  ?, "h�   
  via2  +W� "(   
  via3  -n� �,   
  via3  -&� �,   
  via2  s� 
B�   
  via3  ǜ ��   
  via3  ǜ !   
  via2  � "�    
  via2  �L �|   
  via3  T� �|   
  via4  T� T   
  via2  � �    
  via3  �� �    
  via3  �� !.$   
  via2  ,X ̠   
  via2  �H �   
  via   , 
�,   
  via2  .� 'T   
  via3  "�T 'T   
  via3  "�T !�   
  via3  � Hd   
  via3  �     
  via3  � ""H   
  via2   $� =`   
  via2   � 	�d   
  via3  %�� 	�d   
  via2   j� EP   
  via    j� �x   
  via2  !2 ]T   
  via2  !0 J|   
  via3  "� J|   
  via3  "� ��   
  via2  h @H   
  via3  b� @H   
  via3  b� "Ep   
  via3  -j� �   
  via3  �8 #$   
  via3  �8 "(   
  via2  .Y< ��   
  via2  �� Ԙ   
  via3  #�D Ԙ   
  via3  &�L 
 �   
  via3  &�L �h   
  via2  �( ��   
  via3  �� ��   
  via3  ��  ��   
  via3  U�  ��   
  via3  U� $'�   
  via2  �� )h   
  via3  WP `   
  via2  , $�p   
  via4  	 � $݀   
  via4  #D $݀   
  via3  &�� \   
  via3   Ơ 	�T   
  via3   Ơ EP   
  via2  ��  ��   
  via3  
�h �   
  via2  �  �X   
  via3  S� �X   
  via3  S� @   
  via2   �� )h   
  via2  Y� ��   
  via2  ȼ �l   
  via3  :( �l   
  via3  :( �8   
  via3  Y� �8   
  via4  *�, Y�   
  via3  -d ��   
  via   !�, ��   
  via2  !�, 
 �   
  via3  %0 �   
  via3  -�d m�   
  via3  '�, B�   
  via2  4( !T   
  via3  WP !T   
  via3  WP )h   
  via   $f\ ��   
  via3  ,Ҝ �x   
  via2  ^  Ը   
  via2   o�   
  via3  "� �   
  via   %s� �   
  via2  � �,   
  via3  ˈ �,   
  via2  � #۰   
  via4  *a� b|   
  via2  %�@ ��   
  via3  �x %�   
  via2  &� �   
  via2  #l �p   
  via2  �p  �l   
  via2  �p ]T   
  via3  �H ]T   
  via3  �H ؀   
  via2  � j�   
  via2  +< ]T   
  via3  8 ]T   
  via3  �� B�   
  via3  'T B�   
  via3  'T L�   
  via3  �l ��   
  via3  �l �   
  via2  $ �   
  via4  
� ct   
  via4  
� $�   
  via4  � $�   
  via3  � Y�   
  via3  )�4  �   
  via2  )��  �   
  via4  *4� ��   
  via2  )�� el   
  via3  )�� el   
  via4  )�� �t   
  via4  *# �t   
  via4  *# b|   
  via2  �4 6�   
  via   �l �   
  via4  	N� &�x   
  via2  �� >0   
  via2  �  !C�   
  via3  �� !C�   
  via3  �� "h�   
  via2  �� B�   
  via2  
90 !�(   
  via2  X$  ��   
  via2  *@h %�8   
  via4  �h j�   
  via3  �h �   
  via2  �� �   
  via2  !�$ ��   
  via3  'VP �p   
  via3  �8 ��   
  via2  ݈  �   
  via3  D  �   
  via3  D sX   
  via2  � sX   
  via2  � ��   
  via2   l� ��   
  via3  h� ip   
  via4  h� &�x   
  via2  �� ��   
  via3  �� ��   
  via3  �� ""H   
  via3  $�� j�   
  via3   ~\ �D   
  via2  	5l h|   
  via3  	�H Al   
  via3  �� �   
  via3  	�H Z   
  via3  	�� ��   
  via2  �  ��   
  via   I�  @   
  via2  "�| j�   
  via3  $N� :,   
  via3  |� %�    
  via2  �H �   
  via3  *� �   
  via3  *� #��   
  via4  ,�� -P   
  via2   �X �p   
  via2  �0 $I   
  via2  �0 $%�   
  via4  *� ��   
  via2  #�� ��   
  via3  #"$ ��   
  via3  #"$ �   
  via3  �  [X   
  via2  �� �   
  via2   G� dH   
  via2  _� 9�   
  via2  &�4 ��   
  via3  _� ��   
  via2  � %�(   
  via2  �H !   
  via3  � !   
  via3  wh %�(   
  via4  wh &T�   
  via4  � &T�   
  via3  � &-p   
  via2  �( �   
  via3  O� �   
  via3  O� ��   
  via2  �� �0   
  via2  �X ip   
  via2   I� ip   
  via2   I� ��   
  via2  L cp   
  via3  	�� �p   
  via3  
� $l8   
  via3  
� $I   
  via2  %� %�   
  via2  � B�   
  via2   4$ ��   
  via2  !�� ��   
  via2  )6� ��   
  via3  !� ��   
  via2  #  �    
  via2  � -P   
  via3  ", -P   
  via3  ", Ј   
  via4  *� @�   
  via3   8 	�T   
  via2   � 	�T   
  via2   � ��   
  via2  T@ %�(   
  via2  � �   
  via3  )� �   
  via4  )� ȸ   
  via4  �\ ȸ   
  via3  �\ ��   
  via2  � ��   
  via2  � Ј   
  via4  � &�x   
  via2  � ��   
  via2  	n `   
  via2  
�� �D   
  via3  	)� �D   
  via2  $A@ ��   
  via3  0� ��   
  via2  /H cp   
  via2  !� h|   
  via   !� b|   
  via2  %�� -   
  via3  %�� ]T   
  via2  {� ��   
  via2  �d hx   
  via3  !�H hx   
  via3  !�H �0   
  via4  0� �   
  via   "�� $   
  via   +� $   
  via2  ~� �x   
  via2  8� ��   
  via2  b� �x   
  via2  � �x   
  via   f� "�8   
  via2  #t, up   
  via3  #ht ��   
  via3  #ht Ј   
  via3  #�T Ј   
  via4  #�T &�x   
  via2  !�  �   
  via2  "=� �D   
  via3  %�< �D   
  via3  %�< ��   
  via3  &L� !T   
  via2  �0  �l   
  via2  �l �|   
  via3  !r� �|   
  via3  !r� h|   
  via3  #t, g8   
  via2  �� ��   
  via4  �� ��   
  via3  �� !�(   
  via3  �� �x   
  via3  ��  �   
  via2  ${� `�   
  via3  's� `�   
  via3  's� g�   
  via2  �h j�   
  via3  n� j�   
  via3  n� ��   
  via2  �L ؀   
  via   �� aX   
  via   f� aX   
  via3  (]� �0   
  via2  "߼ �8   
  via2  #/� 	E   
  via3  #� 	E   
  via2  !A� j�   
  via3  "�� j�   
  via3  "�� ��   
  via2  p 8   
  via   �0    
  via2  �8  �l   
  via2  � U�   
  via3  @� U�   
  via3  @� �   
  via2  &^D ��   
  via3  #t, ��   
  via3   ;� ��   
  via4  -i  �   
  via4  .Ox �   
  via3  .Ox ��   
  via2  .,P ��   
  via   .,P R�   
  via2  *�  �\   
  via2  6� �   
  via3  ct �   
  via4  ct ��   
  via4  @L ��   
  via3  @L �   
  via2  s �   
  via   s ��   
  via4  0� k    
  via3  &�H �0   
  via3  %�L ��   
  via3  *�\ 9�   
  via2  &�l �8   
  via4  *W� '   
  via4  *W� J4   
  via4  $  J4   
  via   #�� �x   
  via2  #�� f   
  via3  $;d f   
  via2  3� �   
  via3  `� 9�   
  via3  `� ��   
  via2  � �   
  via2  %Ѥ ��   
  via2  )� o�   
  via2  )� `   
  via3  +� `   
  via3  +� �   
  via2  ,X P0   
  via2  � �t   
  via2  !�p �t   
  via   !�p �x   
  via2  �, "`   
  via2  l@ ��   
  via3  p� ��   
  via3  p�  ��   
  via2  � #۰   
  via3  �, $p    
  via   &�H <d   
  via3  r� ��   
  via3  r� ��   
  via2  	3x �   
  via   	� Z�   
  via   �p Z�   
  via   �p 
�,   
  via   �� ��   
  via2  � Ը   
  via3  �8 Ը   
  via4  �8 &�x   
  via4  �� &�x   
  via2  @ !C�   
  via   �P  @   
  via4  ,0� T`   
  via3  ,0� ̠   
  via3  �< f   
  via4  �< �(   
  via4  !� �(   
  via3  !� f   
  via2  !�D f   
  via2  !�D @   
  via2  �� ��   
  via2  v� �|   
  via3  �� �|   
  via3  �� 8   
  via2  -�� P|   
  via2  � ��   
  via3  RL |�   
  via   4 "�8   
  via2  � ��   
  via   �h  @   
  via2  Rl 	�<   
  via2  Z< |�   
  via3  � |�   
  via3  � ��   
  via2  )�� ��   
  via2  &74 6�   
  via3  '�, 6�   
  via2  R  ��   
  via2  �� "��   
  via2  t !�8   
  via2  �� ��   
  via3  �h ��   
  via3  �h �h   
  via2  �@ f   
  via3  �T "(   
  via4  �T I8   
  via4  N I8   
  via3  N ��   
  via2  &�H �0   
  via   *�� 
�,   
  via   &�l 
�,   
  via   &�l <d   
  via2  � �x   
  via   %�L e    
  via   �X e    
  via2  �� !f�   
  via3  , "��   
  via   �H ��   
  via   �h ��   
  via2  3 �(   
  via3  �, �(   
  via3  �,  ��   
  via2  H !�   
  via   �d  ʈ   
  via2  &@� �x   
  via2  $f\ f   
  via3  %dD f   
  via2  \x t�   
  via2  \x �   
  via2    9�   
  via3  a� 9�   
  via3  a� 8   
  via2  YD EP   
  via2  *@ "(   
  via   �P �x   
  via2  %w� Θ   
  via2  4� Y�   
  via2  %�� �,   
  via3  &L� �,   
  via3  *4� o   
  via2  �� k�   
  via3  � k�   
  via4  � ��   
  via2  YD 	l   
  via3  � 	l   
  via3  � j�   
  via2  ,��    
  via2  *� �8   
  via3  +�� �8   
  via4  -� w@   
  via2  �� ��   
  via2  P �    
  via2  
� �    
  via   
� �   
  via2  �@ \   
  via2  � �   
  via3  
�� �   
  via3  
�� 
B�   
  via2  U ��   
  via4  �� ��   
  via3  �� �p   
  via2  J �    
  via   e� e    
  via   �P e    
  via3  %=4 �   
  via3  %=4 ��   
  via3  G  $�`   
  via2  � ��   
  via2  !f� �h   
  via3  "($ ~�   
  via4  "($ ��   
  via4  -< ��   
  via3  -< Ј   
  via2  A� ��   
  via3  �� ��   
  via3  �� @H   
  via2  �� ��   
  via2  P� H�   
  via3  -� H�   
  via2  G� 9�   
  via2  n� C�   
  via3  �� C�   
  via2  
�( 6�   
  via2  %�� ��   
  via3  %< ��   
  via3  %< Θ   
  via3  N� !�(   
  via3  ؤ !��   
  via4  ؤ !Ĉ   
  via2  b� �H   
  via2  j� �    
  via3  ^l �    
  via3  ^l "(   
  via2  %Z� �   
  via3  �$ cp   
  via2  �� ��   
  via2  %�H ��   
  via3  'u� ��   
  via2  "z, o�   
  via4   >� ܈   
  via2  k  @H   
  via   k  ��   
  via2  
#� ��   
  via2  
'� <d   
  via3  	�$ <d   
  via3  	�$ �x   
  via2  &3L �x   
  via2  %� Q�   
  via3  $� Q�   
  via3  �� !f�   
  via2  �� j�   
  via2  
�� "(   
  via3  
m� "(   
  via3  
m� P   
  via2   �$ �|   
  via2  �� �H   
  via3  � �H   
  via3  � B�   
  via3  *�D ��   
  via2  .� Hd   
  via3   � Hd   
  via4   � Y�   
  via2  �P �X   
  via4  �$ T`   
  via2  %\ ��   
  via2  S� sX   
  via3  $ sX   
  via3  $ #۰   
  via2  }� ��   
  via3  	׈ ��   
  via3  	׈ 8   
  via4  ڼ 	!�   
  via2  .4 ��   
  via3  .*\ ��   
  via4  %ϰ ?�   
  via3  "7� ��   
  via2  3 !�(   
  via4  � !?�   
  via4  �� !?�   
  via   Yd $   
  via3  �� 	p   
  via3  �� 	�d   
  via2  $�� 
F�   
  via2  � 8   
  via2  � ��   
  via3  1� ��   
  via3  1� ��   
  via2  %�l ��   
  via2  %s� �,   
  via2   � �,   
  via2   � 6�   
  via2  �� �   
  via3  @p �   
  via3  @p "��   
  via2  �P !��   
  via2  /� ��   
  via2  &�l j    
  via2  ,m �H   
  via3  '!� �H   
  via2  �\ C�   
  via2  
� j�   
  via3  
  j�   
  via4   | ��   
  via2  
�� Y�   
  via3  &X Y�   
  via   � ��   
  via2  Y� ��   
  via2  N@ $p    
  via2  �� $�`   
  via2  @H !�   
  via2  "`�    
  via3  @H    
  via2  *6� !T   
  via3  !�L !T   
  via3  !�L Y�   
  via   2� �\   
  via2  bx ��   
  via2  �� ��   
  via2  �p �   
  via2  � �   
  via2  � P0   
  via2  .d� j�   
  via2  *�, ��   
  via3  -E� ��   
  via3  
� �x   
  via2  � $l8   
  via2  � ̠   
  via2  � "��   
  via2  b� %�   
  via2  �� �   
  via2  8X �   
  via2  8X �h   
  via2  *y '   
  via2  "S !T   
  via2  �� %�(   
  via3  5D %�(   
  via4  5D &1X   
  via4  "x &1X   
  via3  "x &
H   
  via2  ^� k    
  via2  ^� �   
  via2  
� �x   
  via2   8   
  via2  	N� !*<   
  via3  	q� !*<   
  via4  	q� &�x   
  via2  hx 	�,   
  via   hx 
�,   
  via4  0� Ը   
  via2  "�� B�   
  via4  'm� �   
  via4  ,�L �(   
  via3  ,�L P0   
  via2  )6� D|   
  via3  
�|    
  via3  
�T    
  via3  
�T T�   
  via2  �� Al   
  via2  �� =`   
  via2  �0 ��   
  via2  � ��   
  via3  ~� ��   
  via3  ~� >   
  via2  � >   
  via2  � ��   
  via2  S  �`   
  via2  �� `   
  via3  �t `   
  via3  �t k    
  via3  >� #۰   
  via2  �� !QL   
  via3  4� !QL   
  via2  (�� �4   
  via2  '�� B�   
  via3  (�L B�   
  via3  (�L ��   
  via3  '�� �    
  via3  &�h k    
  via3  &�h �0   
  via3  0� �0   
  via3  &ɰ  �   
  via3  &��  �   
  via2  %h, �   
  via2  r� Y�   
  via   	�$ ��   
  via2  �� ��   
  via2  84 :,   
  via3  z� :,   
  via4  z�    
  via2  $;d 2�   
  via2  
�� 8   
  via3  30 8   
  via4  30 _$   
  via4  �, _$   
  via3  �, 8   
  via2  �$ ��   
  via2  �� �   
  via3  ]t �   
  via3  ]t ��   
  via4  $�$ @�   
  via2  1� �   
  via2  �� "��   
  via   ~@ b|   
  via2  � 	��   
  via2  � �x   
  via2  � H�   
  via3  {� H�   
  via4  {� p    
  via4  �$ p    
  via3  �$ )h   
  via2  ` g�   
  via3  	�� �   
  via3  	�� �   
  via2  	�$ �   
  via4  	�� &�x   
  via2  �� Ј   
  via3  $� Ј   
  via4  $� ��   
  via4  m� ��   
  via3  m� ̠   
  via2  [� @H   
  via2  _� �   
  via3  �� �   
  via4  ��     
  via4  $�4     
  via3  $�4 gX   
  via3  *� ��   
  via2  "� g�   
  via3  $�$ g�   
  via2  'c� ��   
  via3  'm� ��   
  via3  . D4   
  via3  �� #$   
  via4  �� ��   
  via2  �� 	�,   
  via    \ $   
  via2  �� �l   
  via2  �  =`   
  via3  �� =`   
  via3  �� �   
  via2  ,��    
  via2  ,δ �T   
  via3  -�d �T   
  via3  0� �p   
  via3  %Ѥ �D   
  via2  �� 	�,   
  via2  �< �   
  via2  .[0 ��   
  via3  $�0 @H   
  via3  $�0 ��   
  via3  �8 �x   
  via2  �� ��   
  via2  T ~�   
  via2  ~� ��   
  via2  5D �0   
  via3   �0   
  via3      
  via2  $#� ��   
  via2  %H� ��   
  via3  %�� �   
  via3  &-p �   
  via2  �� EP   
  via2  ~ �    
  via2  $� �h   
  via2  (� f   
  via3  .*\ �   
  via3  -�H �   
  via4  0� =8   
  via2  �p %�8   
  via2   � $�`   
  via2  w <   
  via3   <   
  via   ,�D ��   
  via2  & � �D   
  via2  �� �X   
  via3  $� �X   
  via3  $� ��   
  via2  
F� �   
  via   
J� $   
  via2  < �   
  via3  �P �   
  via3  �P ��   
  via2  �H �   
  via2  V4 L�   
  via2  , M�   
  via3  �D M�   
  via3  �D �    
  via2  $�� �p   
  via3  %�� _l   
  via2  $�� �   
  via3  $�D �   
  via2  !� !�(   
  via3  #"$ !�(   
  via4  #"$ ""H   
  via4  *�� ""H   
  via3  *�� !�8   
  via2  ""H ��   
  via2  "&0 sX   
  via3  $�  sX   
  via3  $�  ��   
  via2  � �x   
  via2  � -P   
  via3  �@ -P   
  via3  �@ @H   
  via2  *� ��   
  via2  *� B�   
  via3  *0� B�   
  via2  Wp 5�   
  via2  [X dp   
  via3    dp   
  via2  &� �8   
  via2  �\ #۰   
  via2  M  �   
  via2  &� @H   
  via2  ,i$ ��   
  via2  �� 	�,   
  via3  ׄ 	�   
  via3  ׄ D   
  via2  $�D �   
  via3  � &-p   
  via2  5� ��   
  via2  =� 	�<   
  via2   � RH   
  via2  %�� RH   
  via2  %�� ��   
  via2  )� �   
  via2  )�L EP   
  via3  )X EP   
  via2  �\ !T   
  via2  �\ ؀   
  via3  y\ ؀   
  via3  y\ ��   
  via2  �� ��   
  via   �� ��   
  via3  #=| �l   
  via2  � x�   
  via3  /  x�   
  via4  /  ��   
  via4  "� ��   
  via3  "� x�   
  via2  4 �   
  via3  &X Al   
  via3  &X ��   
  via2  	�� j�   
  via2  	5l �8   
  via2  Q &-p   
  via3  Z� &-p   
  via4  Z� %�   
  via4  � %�   
  via3  v� @H   
  via4  v� gX   
  via4  &L� gX   
  via3  &L� @H   
  via2  J  �   
  via3  �L  �l   
  via3  �L ]   
  via2  nx @H   
  via2  r` gX   
  via3  t gX   
  via4  t @H   
  via4  ]� @H   
  via3  ]� gX   
  via2  !�l ��   
  via3  #=| ��   
  via2  �� �x   
  via2  �    
  via2  *�x )h   
  via3  *� ��   
  via2  *�p ��   
  via2  #�� Θ   
  via   $N� 
�,   
  via2  �  �\   
  via3  �  �\   
  via3  � �D   
  via2  �� �   
  via2  ո ��   
  via3  �L ��   
  via3  �L aX   
  via2  �� @H   
  via3  ., �x   
  via3  ., gX   
  via2   gX   
  via    aX   
  via2  $T �0   
  via2  #` RH   
  via2  !G� �   
  via2  �� o�   
  via2  -� ��   
  via2  -�  P|   
  via2  -G� ��   
  via2  -"� @H   
  via2  �T �x   
  via2  � �   
  via3  �8 �   
  via3  $�  �p   
  via2  �� ��   
  via2  � ��   
  via2  "�� ��   
  via2  "�� �l   
  via2  ]� =`   
  via3  :� ��   
  via2  0� ��   
  via2  +d -   
  via2  *�l EP   
  via3  +	� EP   
  via2  #G@ 8   
  via2  "h� f   
  via2  9� -   
  via2  SH �x   
  via3  �< <   
  via2  	)� <   
  via2  	)� `   
  via2  *� j�   
  via2  #�� D|   
  via2  � �h   
  via3  �\ �h   
  via3  �\ )h   
  via2  cp 	l   
  via   ed $   
  via2  �t ��   
  via3  �� `�   
  via2  &�� _l   
  via2  $�� ��   
  via3  $�  ��   
  via2  @ �4   
  via2  �D �4   
  via2  �D ��   
  via2  �l ��   
  via2  �l 
�D   
  via2  �d 
�D   
  via   �d ��   
  via3  RL �l   
  via2  y8 !T   
  via2  �p !T   
  via   �p $   
  via2  �, +<   
  via3   � 'T   
  via4   � Nd   
  via4  �< Nd   
  via2  >� T�   
  via2  
�� =`   
  via3  >� =`   
  via3  >� FL   
  via3  |� 
�l   
  via2  |� �   
  via2  k� "A�   
  via2    !f�   
  via2  � �0   
  via2  �d h�   
  via3  �< h�   
  via2  � �h   
  via3  0 �h   
  via3  0 �   
  via3  � ��   
  via2  �� �   
  via2  C� aX   
  via2  j$ ��   
  via2  (#d �   
  via2  &� ��   
  via2  , �   
  via2  R  !��   
  via2  "� ��   
  via2  �� up   
  via2   zt 
�d   
  via2  !�t 6�   
  via3  $�� 6�   
  via2  v &
H   
  via2  �@ !�8   
  via2  � $%�   
  via2  MH �   
  via2  L 	��   
  via3  I� 	��   
  via2  �L D   
  via2  � �0   
  via2  -,t ��   
  via3  �� !�(   
  via3   >� @H   
  via2  #l %�   
  via2  Rl �8   
  via3  �x �8   
  via2  
8  �   
  via2  Nd  �   
  via2  Nd �   
  via2  �  �x   
  via2  j$ 
 �   
  via2  .Ql �X   
  via2  ,�\ �p   
  via3  *� �p   
  via3  *� ��   
  via2  ,�4 Θ   
  via2  	N� >0   
  via2  ~� ~�   
  via2  G  �   
  via2  �� sX   
  via2  �X 
�   
  via2  }� ��   
  via3  �0 ��   
  via4  �0 9�   
  via4  @L 9�   
  via2  \ ��   
  via2  D !T   
  via2  Z� ��   
  via2  �� D|   
  via2  
p �   
  via2  �� !�8   
  via3  �� !�8   
  via4  �� &�x   
  via   W� ��   
  via   "� �\   
  via2  �, !�(   
  via2  
� !�   
  via3  	)� <   
  via2  .d� $L�   
  via2  T� �   
  via2  %� "�    
  via3  �� "�    
  via4  �� # 0   
  via4  �� # 0   
  via2  �P 	l   
  via2  �8 
B�   
  via2  �< )h   
  via2  �H FH   
  via3  �  FH   
  via2  �( #۰   
  via2   $L�   
  via2  o� ��   
  via2  � ��   
  via2  *<� ��   
  via2  *DP ��   
  via2  � Y�   
  via2  d 
f   
  via3  W 
f   
  via3  � �    
  via2  �x %�   
  via4  � �   
  via3  
� dp   
  via2  `� dp   
  via2  `� 	�T   
  via2  �� 8   
  via2  H �|   
  via2  �t ��   
  via2  �� ��   
  via2  �� �`   
  via2  �� "��   
  via2  "� [X   
  via2   G� �@   
  via3  "� �@   
  via3  "� )h   
  via2  �� �   
  via2  �� Y�   
  via3  $^� :,   
  via3  w &�x   
  via2   <   
  via2  �� ��   
  via2  �| �   
  via2  #z o�   
  via2  )>� 6�   
  via3  *� 6�   
  via3  *� j�   
  via   _d $   
  via2  
�P 	h4   
  via4  	� 	A$   
  via3  	� 	�T   
  via2  �d 	�T   
  via   �d ��   
  via2  
� $%�   
  via2  � EP   
  via3  �� EP   
  via3  �� �x   
  via2  C� 6�   
  via2  C� it   
  via3   | it   
  via2  `� �X   
  via   ň ��   
  via3  
!� �   
  via2  �� `�   
  via2  �� �,   
  via4   4� &0   
  via3  	 � !�   
  via3  	 � $�p   
  via2  x #$   
  via2  U\ g�   
  via2  > 	l   
  via2  
H� 9�   
  via3  
�� 9�   
  via4  
�� �   
  via2  �� 	l   
  via2  ֬ ��   
  via2  _d ��   
  via   �  b|   
  via   
ɸ b|   
  via2  e� �(   
  via2  6� |�   
  via2  ]t |�   
  via2  ]t �h   
  via2  �p ��   
  via2  ܬ 6�   
  via3  �� 6�   
  via4  �� |   
  via4  #� |   
  via3  #�  �l   
  via2  �� Al   
  via2  �X ��   
  via3  
!� ��   
  via2  
� j�   
  via2  p hx   
  via2  �  \   
  via2  !
� 
F�   
  via2  *�D ��   
  via2  )�| Y�   
  via3  *�D Y�   
  via2  �( �(   
  via4  ,Ҝ ��   
  via2  �d �0   
  via3  ,� �0   
  via3  ,� �8   
  via2  $�� 
#�   
  via3  $� _l   
  via2  7� =`   
  via2  QP �p   
  via2  � ɔ   
  via2  �� !�   
  via3  �\ !�0   
  via4  �\ !�   
  via4  �d !�   
  via3  �d !��   
  via2  &�  ��   
  via2  ''p 	�|   
  via2  �� j�   
  via2  � #$   
  via2  +� #$   
  via2  +� �X   
  via2  )�p ��   
  via2  )� �|   
  via2  �� �0   
  via2  �� �0   
  via2  Q ��   
  via2  � �0   
  via   �$ �x   
  via   f� �x   
  via2  f� �   
  via2  �$ ��   
  via3  �� ��   
  via3  �� ��   
  via2  6D @H   
  via2  �� ��   
  via3  �� ��   
  via2   � !�(   
  via2  #�� !��   
  via2  
 �h   
  via2  �$ �   
  via4  #EL &^D   
  via2  )�� &74   
  via2  8� �|   
  via2  �H  {   
  via3  ��  {   
  via3  �� x�   
  via2  ;� x�   
  via2  ;� ��   
  via2  	�t !�   
  via3  x@ &
H   
  via4  x@ &1X   
  via4   4� &1X   
  via2  �� �   
  via3  .� Al   
  via4  �$ �   
  via2  E, �   
  via3  � �   
  via3  � �   
  via    �  b|   
  via2  #� ��   
  via2  V0 �   
  via2  +:h �x   
  via2  ,6\ o�   
  via2  %� "��   
  via2  #?p "��   
  via2  �$ `�   
  via3  �l ��   
  via2  ,�D j�   
  via2  !�$ !T   
  via2  !�$ ��   
  via2  )%4 �@   
  via2  (%X �   
  via3  (�� �   
  via2  s\ Hd   
  via2  
Zd ��   
  via3  � ��   
  via2  Q !�8   
  via2  �| <�   
  via2  &͘ 
%�   
  via2  '�H \   
  via3  ) \   
  via4  ) jp   
  via4  .� jp   
  via2  M  !*<   
  via3  ݬ !*<   
  via3  ݬ #۰   
  via2  o 	l   
  via2  
y� ��   
  via2  
V| ��   
  via   
V| 
�,   
  via2  #`� �   
  via2  |� `�   
  via3  �� `�   
  via4  �� ��   
  via4  |� ��   
  via2  %�H ��   
  via   !� �(   
  via2  !h� !T   
  via2  �@ �|   
  via2  �� �0   
  via2  9� ��   
  via2    ��   
  via2  !�� �   
  via2  h� �   
  via   V� <d   
  via   �$ <d   
  via2  �$ j�   
  via2  @p �H   
  via2  6� H�   
  via2  5� -   
  via2  �� �,   
  via3  | �,   
  via2  �\ $�   
  via2  �d  �l   
  via2  �d  �4   
  via3  &�  �4   
  via3  &�  �   
  via4  ,4h ɔ   
  via2  , `   
  via3  ,p� `   
  via3  ,p� j�   
  via2  
7< 	!�   
  via2  �� K0   
  via3  Y� K0   
  via4  Y� �   
  via4  !x �   
  via3  !x �   
  via2  �@ �   
  via3  ]� ��   
  via4  ]� ��   
  via4  !Ĉ ��   
  via3  !Ĉ ��   
  via2  �  �l   
  via2  �� z|   
  via2  "
� ��   
  via2  LH A�   
  via3  � A�   
  via2  � 9�   
  via2  Ș ]T   
  via2  :� ��   
  via2  �� ��   
  via2  � ׬   
  via2  ��  �l   
  via2  5$ �    
  via2  	�  6�   
  via3  �� 6�   
  via4  �� kD   
  via4  . kD   
  via2   �� �X   
  via2  �d �X   
  via2  �d �@   
  via3  �� �@   
  via3  �� @   
  via2  (3 ��   
  via2  )uH o�   
  via3  
 � ��   
  via2  � $)�   
  via2  � ��   
  via2  +�� @   
  via2  +v� =�   
  via3  +�� =�   
  via2   �� ��   
  via2  !	 el   
  via2  *DP ��   
  via2  $ی �   
  via2  e  
B�   
  via2  v( 
�   
  via2  *�� ��   
  via2  �( ��   
  via2  �� ��   
  via2   M� 
�l   
  via2  jp #۰   
  via2  � !QL   
  via2  n0 �H   
  via2  �      
  via2  �� �H   
  via2  � &
H   
  via2  "� !�8   
  via3  E� !�8   
  via3  | -   
  via2  �� �H   
  via2  � ��   
  via4  'u� ��   
  via2  �� [X   
  via2  �  "`   
  via3  � $٘   
  via3  �, $٘   
  via3  �, &
H   
  via2  �� &-p   
  via2  �� %�8   
  via2  -�8 	l   
  via2  ,�� )l   
  via3  -�� )l   
  via   -�� ��   
  via2  ��  �<   
  via2  �D  ,�   
  via3  `�  ,�   
  via4  `�  S�   
  via4  Ѩ  S�   
  via2   ��   
  via2  kD gX   
  via2  �� �   
  via2  n0 �   
  via2  �< �   
  via2  � ��   
  via3  � ��   
  via3  � k    
  via2  "�0 �p   
  via3  "7� �p   
  via2  ,M� �   
  via2  +z� 8   
  via2  e� ��   
  via2  84 ��   
  via2  �$ &-p   
  via3  ,| &-p   
  via4  ,| &`   
  via4  �� &`   
  via3  �� &-p   
  via4  �d #$   
  via4  �P #$   
  via2  #-� j�   
  via2  #Q EP   
  via2  �l �d   
  via3  < �d   
  via3  < 	�,   
  via2  � 	�,   
  via   � ��   
  via2  m� -   
  via2  	p %�   
  via3  	�� %�   
  via3  	�� Px   
  via2  %X� "d�   
  via2  #� "A�   
  via2  �� 	E   
  via2  �� 
B�   
  via2  � 
B�   
  via2  � �   
  via2  �� A�   
  via2  �p #$   
  via3  ^H #$   
  via2  q� �d   
  via2  F� ��   
  via3  q� ��   
  via2  ?, :,   
  via3  O :,   
  via3  O `�   
  via2  oP �   
  via3  �d �   
  via2  �� �   
  via2  �� ��   
  via3  � ��   
  via4  � ��   
  via4  GD ��   
  via3  GD #$   
  via2  $ #$   
  via2  $ �   
  via2  	f@ �(   
  via3  	p �(   
  via4  	p �8   
  via4  Q� �8   
  via3  Q� �(   
  via2  .� �(   
  via2  .� D   
  via3  �� 	�|   
  via2  �� 	�|   
  via   �� 
�,   
  via2  ��    
  via2  � �   
  via2  �� �   
  via2  ո :p   
  via2  ', o�   
  via3  � o�   
  via3  � FL   
  via2  R� �   
  via3  �( 9�   
  via2  "/� ��   
  via   "/� ]�   
  via2  :� �l   
  via2  � �X   
  via2  �L 9�   
  via3  =� 9�   
  via3  =� dp   
  via2  '0 �x   
  via2  'D� ��   
  via2  "�� D   
  via   ", �(   
  via3  E� &0   
  via2  u %�(   
  via3  O� %�(   
  via3  O� &-p   
  via2  � 8   
  via2  U 8   
  via3  �� 8   
  via2  c �x   
  via2  )sT $L�   
  via2  Ԝ k    
  via3  �� k    
  via3  �� �   
  via2  |� �   
  via   |� ��   
  via  �  B�        .� &�\ +  ,VR_NO_BUS    
  via2  vp �   
  via2  � �   
  via2  � -   
  via2  
N� Y�   
  via2  
N� ��   
  via3  �X Px   
  via2  �� �X   
  via   !�� ��   
  via2  (�� �\   
  via2  )y0 j�   
  via2  �| d�   
  via2  Z@ �   
  via3    �   
  via3    cp   
  via4  0� ̠   
  via3  (��    
  via3  (�� ��   
  via2  C� j�   
  via2  &\ ��   
  via2  �L ��   
  via   �L ��   
  via   c ��   
  via2  +B8 !�(   
  via   +@  ʈ   
  via2  !�, \   
  via2  !�� 
j   
  via3  �X @H   
  via2  4 Px   
  via2  �X Ҁ   
  via2  �� �p   
  via2  \4 �x   
  via2  \ P   
  via2  b %�   
  via2  kh �H   
  via2  "�� `�   
  via2  "� �D   
  via2  !�� �D   
  via3  _� 9�   
  via2  �� �P   
  via3  5� �P   
  via3  5� ��   
  via2  �, Y�   
  via2  $� ��   
  via2  � 
�D   
  via2  �h 
�   
  via3  
 � 
�   
  via2  �H �D   
  via   bT 0D   
  via2  �x 	l   
  via3  &� 	l   
  via2  Ș ��   
  via2  ̀ aX   
  via2  Yh �   
  via3  � �   
  via3  � 	l   
  via2  8� j�   
  via3  *# ��   
  via3  *#    
  via2  '�� o�   
  via2  '�� EP   
  via2  Z� gX   
  via2  -� k@   
  via2  -� !�8   
  via2  �t 8   
  via2  �� Ը   
  via2  �$ Ը   
  via   �$  ʈ   
  via3  DT 6�   
  via3  DT ��   
  via2  !, ��   
  via   !, ��   
  via3  )�� ��   
  via3  �, �   
  via3  �, j�   
  via2  �� �h   
  via   �� '   
  via2  � j�   
  via2  � "p   
  via2  ֬ ��   
  via2  �x j    
  via3  � j    
  via2  � 
f   
  via4  &�� ��   
  via3  &�� ʴ   
  via2  &� ʴ   
  via2  &� ��   
  via2  x� |   
  via2  [� Y�   
  via2  �0 %�8   
  via2  L$ "`   
  via3  D "`   
  via3  D $��   
  via3  � "��   
  via3  #�D @H   
  via2  *�� �h   
  via2  %�� ��   
  via2  oL 6�   
  via3  *� Θ   
  via2  +� `�   
  via2  7� ��   
  via2  �� ��   
  via   �� e    
  via2  -j� `�   
  via2  %�D �T   
  via2  -j� ��   
  via2  -G� ��   
  via2  -G� ��   
  via2  � �   
  via2  � |�   
  via2  !] 5�   
  via3  !�� 9�   
  via4  !�� ��   
  via   $/� �`   
  via2  $?L �8   
  via2  �� �0   
  via3  �, �   
  via3  �, s�   
  via2  %� !�(   
  via2  ({H �   
  via2  �, #$   
  via3  �, #$   
  via3  �, FL   
  via3   | FL   
  via2  �� D   
  via2  !� |�   
  via2  "� T   
  via3  *� D   
  via4  *e� �,   
  via3  *e� �<   
  via2  *�, �<   
  via2  *�, h|   
  via2  �4 �d   
  via2  �� :,   
  via2  x� ��   
  via2  �� g�   
  via2  ְ j�   
  via2  Y� j�   
  via2  Y� ��   
  via2  #�8 #۰   
  via2   �� "�    
  via2  q� `�   
  via2  �d �l   
  via2  '� A�   
  via   -� ��   
  via2  
� 
F�   
  via2  �� !�(   
  via2  #H "`   
  via2   �� $݀   
  via2   � $��   
  via2  $� ��   
  via3  $�� �   
  via4  $��    
  via4  )<�    
  via3  )<� �   
  via2  &� Al   
  via3  &0 Al   
  via4  &0 �,   
  via2  !� wD   
  via3  $�� 
�d   
  via4  $�� 
�t   
  via4   �� 
�t   
  via3   �� 
�d   
  via2  i, &
H   
  via2  	E %u�   
  via3  j� �   
  via3  ְ 	�,   
  via3  ְ 
B�   
  via3  N 
B�   
  via2  �` ��   
  via2   ��   
  via2  �( 
�D   
  via2  � �   
  via3  � %    
  via   !� ��   
  via2  ? |�   
  via2  MH  �\   
  via2  U U�   
  via2  .4 )l   
  via3  &; ��   
  via2  �� \   
  via2  7� �T   
  via2  d ��   
  via2  � =`   
  via2  -	L ��   
  via2  �� �0   
  via3  �d �0   
  via3  �d ��   
  via2  !`� %�(   
  via2  $� $�p   
  via3   �P $�p   
  via2  �L �   
  via2  $� �   
  via2  '� �   
  via2  2� �D   
  via2  �t o�   
  via2  `� 2�   
  via2  ޤ C�   
  via2  	� ��   
  via2  ^� %    
  via3  f` %    
  via4  f` %C   
  via4  � %C   
  via2  ^l |   
  via2  �@ �D   
  via2  �     
  via2  )l Hd   
  via3  �� "��   
  via2  E� �0   
  via2  'q� !�(   
  via2  $   �   
  via2  "�  �l   
  via3  #�  �l   
  via4  #�  ,�   
  via4  '��  ,�   
  via3  '��  S�   
  via2  � �h   
  via    � aX   
  via2  � _@   
  via2  	\ "(   
  via2  	� �   
  via3  
`@ �   
  via4  
`@ J4   
  via4  �( J4   
  via3  �( #$   
  via2  � @   
  via2  �\ "��   
  via3  " "��   
  via4  " "�   
  via4  	5l "�   
  via3  	5l "��   
  via2  	�� "��   
  via2  	�� #۰   
  via2  � �   
  via2  �� �D   
  via2  �� #۰   
  via2   � #H   
  via2  �T 
�l   
  via3  l� ��   
  via3  l� =`   
  via2  $^� j�   
  via2  &�0 #۰   
  via2  (�� "d�   
  via2  �L  �l   
  via2  � �   
  via2   x�   
  via2  �� ��   
  via2  �8 �x   
  via3  	ϸ %�    
  via4  	ϸ &�x   
  via2  (RD 	l   
  via2  (V, ��   
  via3  �� $�   
  via2  � $�`   
  via3  �� $�`   
  via4  �� &�x   
  via2  � D|   
  via2  T� L�   
  via2  qh ۔   
  via2  %N� �   
  via2  '5 @   
  via2  ,8P �   
  via3  0� �   
  via3  ut 	�,   
  via   �� 0D   
  via2  �� x�   
  via2  (i� �    
  via2  v 
��   
  via3  
�h 
��   
  via2  %�t 6�   
  via2  � ��   
  via2  �l `�   
  via2  �� "h�   
  via2  #�� ��   
  via2  � #۰   
  via2  �� $�   
  via2  �P �   
  via2  	�� %�    
  via2  +�� )h   
  via3  ,�� �    
  via2  -C� h|   
  via2  (�� �D   
  via2  ,@ �   
  via2   C�   
  via3  � C�   
  via3  � ��   
  via2  6� Al   
  via3  �  ET   
  via3  �  `�   
  via2  S  	E   
  via3  
A  	l   
  via4  
A  	�<   
  via4  ut 	�<   
  via2  ,� ��   
  via2   ;� T   
  via2  ~d ��   
  via2  	�    
  via2  �0  �l   
  via   kd 0D   
  via2   � #۰   
  via2   � $%�   
  via2  �8 �   
  via2  X L�   
  via2  �L �   
  via3  )��  :�   
  via3  )��  :�   
  via2  )P,  �\   
  via2  )W� ��   
  via2  �� ��   
  via2  [� �    
  via2  �  ��   
  via2  7� 
�l   
  via2  �X %�8   
  via2  �@ &�x   
  via2  �0 ��   
  via2  � k�   
  via2  
 �x   
  via3  �� �x   
  via3  �� !tt   
  via2  � Y�   
  via2  �� �H   
  via2  ٠ 	�,   
  via2  	� 
j   
  via2  wd ��   
  via   !, �\   
  via2  �� �h   
  via2  m� %�(   
  via   � $��   
  via2  � !�   
  via2  � "`   
  via2  &ɰ ��   
  via2  ({H 
%�   
  via2  ( D   
  via3  (� D   
  via4  (� ?T   
  via4  ,�L ?T   
  via2  �X #H   
  via2  �0 "��   
  via2  &� �   
  via2  s 
j   
  via3  )�� &\   
  via   �H �    
  via4  : ��   
  via4  : w�   
  via4  �X w�   
  via2  �D l   
  via2  cP ��   
  via3  ,�L D   
  via2  �H Θ   
  via3  [ #$   
  via2  	�  �    
  via2  c� Al   
  via2  -"� ��   
  via2  #�� ��   
  via3  �l `�   
  via2  �� �    
  via2  � 
ϔ   
  via3  �$ ��   
  via4  �$ 
�|   
  via4  �� 
�|   
  via4  �� 
��   
  via4   
��   
  via2  �p D   
  via2  � |�   
  via2  )�4 �   
  via3  %�L �   
  via3  %�L 6�   
  via2  �x �X   
  via2  �� @H   
  via2  Ҁ @H   
  via2  Ҁ gX   
  via2  (sx     
  via2  '�� Θ   
  via2  (+4 �   
  via2  '�\ �   
  via2  ��     
  via2  � �    
  via2  �� |   
  via3  S� |   
  via3  S�  �4   
  via2  &ό !�8   
  via2  #�� "d�   
  via2  #�� ��   
  via2  �� $)�   
  via2  $� �    
  via2  �@ ��   
  via2  $�� 
�d   
  via2   �P wD   
  via2  � !�   
  via2  �� "��   
  via2  �� n0   
  via2  a� l   
  via2  � �,   
  via2  �� :,   
  via2  !� �,   
  via2  !� �   
  via3  %� ��   
  via2  &� 
#�   
  via2  /H ��   
  via2  $ :,   
  via2  (� ��   
  via2  z0 �l   
  via2  �8 `�   
  via2  �� `�   
  via2  &�� ��   
  via2  &o� P0   
  via2  %�� 9�   
  via2  ,� �X   
  via2  �� @   
  via2  #t, ��   
  via2  +�� �   
  via2  )�l ��   
  via2  :, $�H   
  via   � ��   
  via   � ��   
  via2  �x 9�   
  via2  �t  �\   
  via3  p  �\   
  via4  p |   
  via4  ^$ |   
  via3  ^$  �l   
  via2  $�p #۰   
  via2  &
H "��   
  via   )�\ b|   
  via2  $K �    
  via2  $�� j�   
  via2  %Ѥ 
�d   
  via2  �d �   
  via2  G� ��   
  via2  "�� j�   
  via2  (H� L�   
  via2  %�� g�   
  via2  [ 	��   
  via2  r� `�   
  via3  Kt `�   
  via2   ʈ ��   
  via2  '�� f   
  via2  +S� f   
  via2  +S� )h   
  via2  o� D   
  via2  s� >   
  via2  �L  �\   
  via   �� ��   
  via3  �P �   
  via2  ^l 
f   
  via3  %�     
  via3  %� �l   
  via2  �    
  via2  $Ӽ �l   
  via2  +X �   
  via2  �L ��   
  via2  \ l   
  via2   $l8   
  via2  �\ "�    
  via2  ~� �   
  via2  { �|   
  via   �t ��   
  via2  �� ��   
  via2  Xl �   
  via3  R� �   
  via3  R� �   
  via2  '�d &   
  via2  (�� $�   
  via2  &3L %�8   
  via2  'o� #�t   
  via3   &�x   
  via2  "z, �   
  via2  "�� �   
  via2  [X �   
  via2  I� \   
  via2  :� 
j   
  via2  � #$   
  via2  o �   
  via2  ~� ��   
  via2  �8 �   
  via2  	�\ 
��   
  via2  �� H�   
  via2  [� �   
  via2  
`@ @   
  via2  uL �X   
  via   � �x   
  via2  &| 	��   
  via2  �H !.$   
  via2  �\ $l8   
  via2  ] "d�   
  via2  S  !*<   
  via2  �H !*<   
  via2  �H !�8   
  via3  � %�    
  via2  � �x   
  via2  �` ��   
  via2  �D !�(   
  via2  " !�   
  via2  " "h�   
  via2  �� @H   
  via2  )�� �   
  via2  +�$ �|   
  via2  (�X #�t   
  via2  *{  $p    
  via2  
m� "��   
  via4   "��   
  via2  �x �x   
  via2  d aX   
  via4  R� &
H   
  via3  R� %�8   
  via2  GD �0   
  via2  7� �X   
  via2  ! x @H   
  via3   �P P0   
  via2  '� 
�D   
  via3  /� 
�D   
  via3  /� �   
  via2  < 	E   
  via2  @  
ϔ   
  via2  �� 9�   
  via2  MH �4   
  via2  �h #۰   
  via3  � #۰   
  via2   �  J   
  via3   �( J   
  via2  �l �   
  via    ��   
  via2  �� FL   
  via2  �\ ��   
  via2  2\ !�   
  via2  'x �(   
  via2  � ��   
  via2  ژ �l   
  via2  I� �l   
  via2  +�4 Y$   
  via2  �@ $�   
  via3  �t %�8   
  via4  �t &
H   
  via2  �� @H   
  via3  1� @H   
  via3  1� ��   
  via2  !, z|   
  via2  �� ��   
  via2  X� ��   
  via2  �� ��   
  via2  |� o�   
  via3  �d o�   
  via4  �d ��   
  via4  $@ ��   
  via3  $@ ��   
  via2  �� @H   
  via2  k� "A�   
  via2  !�� Ј   
  via3  �� !��   
  via3  �� "`   
  via2  	X ��   
  via2  �P +<   
  via2  $�� 	l   
  via2  �P "`   
  via2  +� �   
  via2  x� n0   
  via2  Al ��   
  via2  rd �   
  via2  � �h   
  via2  	  �x   
  via2  -�� �0   
  via2  $ 	�T   
  via2  �� ��   
  via2  �� 	E   
  via2  � `�   
  via2  l� ��   
  via2  �H 8   
  via2  *L Al   
  via2  (�L Al   
  via2  (�L �   
  via2  �� �d   
  via2  b� �`   
  via2  .M� ��   
  via   -�� ��   
  via2  Td ��   
  via2  w� ��   
  via2  w� :,   
  via2  �@ !�   
  via2  ]� 9�   
  via2  �� ��   
  via2  )_� -   
  via2  (]� ��   
  via3  (�$ ��   
  via2  ('L ��   
  via2  $n, ��   
  via2  %�� ��   
  via2  �4 gX   
  via2  � ��   
  via2  �� "��   
  via2  f` "�    
  via2  g\ ��   
  via2    j�   
  via2  \ >   
  via2  �� Ҁ   
  via2  "�8 �0   
  via2  "�  )h   
  via2  ,� �   
  via2  �, x�   
  via3  J0 Al   
  via2  �\ 	E   
  via2  Q0 !Md   
  via2  ?� "d�   
  via2  z� ��   
  via2  �� l   
  via   �l ��   
  via2  �� �    
  via2  �� j�   
  via2  u( ��   
  via2  
Xp  �l   
  via2  
\X 6�   
  via2  �� ��   
  via2  	� "(   
  via2  � �    
  via2  �, r   
  via3  �� r   
  via3  �� �h   
  via   ct e    
  via2  � ��   
  via2  � ��   
  via2  �H �   
  via2  /� �    
  via2  }� Y�   
  via2  $ � ��   
  via4  YD 
�|   
  via3  YD ��   
  via2  #�d $�   
  via3  "�T $�   
  via3  "�T $I   
  via2  "�D @H   
  via2  #�L �   
  via2  �    
  via2  x� �h   
  via2  *@ EP   
  via2  :( 
�<   
  via2  #`� �   
  via2   �� 2�   
  via2  ,� 
�,   
  via2  �� 	��   
  via2  ,�� �   
  via2  Ȝ `�   
  via4  �, =�   
  via2  �� j�   
  via2  6� �l   
  via3  �4 T�   
  via3  �4 `�   
  via2  �$ ��   
  via2  l� ��   
  via   {P '   
  via2  �x �X   
  via2  F� Al   
  via2  v� ��   
  via3  �� ��   
  via4  �� 
�|   
  via2  6� jp   
  via3  �� jp   
  via3  	�� Z   
  via2  �X AH   
  via2  K� ��   
  via2  D  �   
  via2  -�� r@   
  via2  (�\ D   
  via2  Ll &
H   
  via2  Ր $��   
  via2  � $l8   
  via2  s\     
  via2   @H   
  via2  �\ @H   
  via   �\ �    
  via2  �� ��   
  via2   
f   
  via   �� $   
  via2  P �   
  via2  *S� o   
  via2  *Y� |�   
  via3  *4� |�   
  via2  kd 	!�   
  via3  4 	!�   
  via3  4 ��   
  via2  �� �h   
  via3  � �h   
  via3  � !�(   
  via2   20 �   
  via2   � ��   
  via2  � 	l   
  via2  � 	�,   
  via3  �� 	�,   
  via4  �� 	A$   
  via4  
d( 	A$   
  via3  
d( 	h4   
  via2  !	 ��   
  via2  � o   
  via2  �� C�   
  via2  
�, !�8   
  via2  �� !QL   
  via2  )a� Ј   
  via2  (�� ��   
  via2  
o� �   
  via2  � AH   
  via2  �8 �(   
  via2  �� �4   
  via2  �� 
�,   
  via2  _d ��   
  via2  � 2�   
  via2  � 9�   
  via   �� �   
  via2  > ~�   
  via2  �� ��   
  via   4� �x   
  via2  X �   
  via2  ,�� �h   
  via2  ,��  �   
  via2  �� "(   
  via2  �� aX   
  via2  l� �h   
  via2  )�4 ��   
  via2  ,o  \   
  via2  	�\ ʴ   
  via2  � ��   
  via2  � ��   
  via2  *� C�   
  via   �� e    
  via2  ,�t @H   
  via3  +� @H   
  via3  +� �x   
  via2  << T�   
  via3  � T�   
  via3  � ��   
  via2  	�$ ��   
  via3  � :,   
  via3  �    
  via2  f� ��   
  via3  �� ��   
  via3  �� 9�   
  via2  $ ��   
  via2  �d ��   
  via2  ~  �l   
  via2  �  	�   
  via2  	�L �x   
  via2  ň l   
  via2  �  �   
  via2  � �(   
  via2  �0 !��   
  via2  �� D   
  via2  Č D   
  via2  $� D   
  via   $� e    
  via2  %n ��   
  via2  $�� �`   
  via3  %� �`   
  via2  �@ "��   
  via2  )� !�   
  via   )��  ʈ   
  via2  �� %�8   
  via2  � $�`   
  via2  b� ��   
  via2  � -   
  via2  �D |   
  via2  �� :,   
  via2  _� U`   
  via2  �� o�   
  via2  1� o�   
  via3  #� o�   
  via3  #� ��   
  via2  �� 	l   
  via2  �� ��   
  via2  +؜ 	u�   
  via   +cl b|   
  via2  	�� �   
  via2  	h4 �   
  via3  ٠ �   
  via3  ٠ ��   
  via2  !QL 	E   
  via2  	�� Y�   
  via2  d$ �   
  via2  �� 
�<   
  via2  up #۰   
  via2  �L #۰   
  via2  �L $�   
  via2  �4 %�(   
  via2  
�, &P�   
  via   �d    
  via2  �  �l   
  via2  ��  �l   
  via2  �� 2�   
  via2  ~@ 	E   
  via    \ b|   
  via2  ��    
  via2  � `�   
  via2  �X �H   
  via2  �@ �    
  via2  -?� $�   
  via2  )�| &
H   
  via2  \ &
H   
  via2  �� !�   
  via2  -0 9�   
  via2  !0 ��   
  via2  � �    
  via3  2� �    
  via2  �� �   
  via2   � �   
  via2    ��   
  via2  $  �p   
  via2  88 )�   
  via2  !I| ��   
  via2  U� �0   
  via2  [\ "(   
  via2  � l   
  via2  [� H�   
  via2  �p !�(   
  via2  -X ��   
  via2  �d @   
  via2  '� ��   
  via2  -�p �   
  via2  ,�� :p   
  via4  .Y< #��   
  via2  )� $�   
  via2  -G� @   
  via2  '  j    
  via3  '�� �   
  via2  .�t @H   
  via2  j$ @H   
  via2  f< �0   
  via   E� e    
  via2  dH �   
  via2  'e� ��   
  via2  &�, �H   
  via3  'T �H   
  via2  |� @   
  via2  
h �@   
  via2  %T ��   
  via4  � &�x   
  via2  � ��   
  via2  !C� �0   
  via2  D� 	!�   
  via2  {� j�   
  via3  �� j�   
  via3  �� d�   
  via2  %�� #۰   
  via2  "�� #H   
  via2  � �x   
  via2  �� �X   
  via2  
�X �x   
  via2  � 	l   
  via2  RH |   
  via2  $N� �   
  via3  $r �   
  via4  $r 7�   
  via4  '�� 7�   
  via2  �| j�   
  via   *FD    
  via2  *>t �l   
  via3  )�$ �l   
  via3  )�$ h|   
  via2  *L h|   
  via   *L b|   
  via2  |� �   
  via3  -�H )l   
  via2  �� L�   
  via2  �$ @H   
  via2   ��   
  via2  @ �d   
  via2  1� 
j   
  via2  � ��   
  via2  �H ��   
  via2  �� �0   
  via2  �L h|   
  via2  ϴ �   
  via2  � �h   
  via2  �4 ��   
  via2  �� ��   
  via2  	%� ��   
  via2  	%� ��   
  via2  'o� Al   
  via2  "� ��   
  via2  !T �0   
  via2  � P   
  via2  7� �   
  via2  �| k    
  via2  �D ��   
  via2  �l 	�,   
  via2  )�     
  via2  +Q� �   
  via2  +s �    
  via2  +(� D   
  via2  )� �    
  via2  �� �0   
  via2  � �X   
  via2  �` aX   
  via2  $� @H   
  via2  C� s�   
  via2  %�� �   
  via3  �� ��   
  via2  �\     
  via2  �< �d   
  via3  �d �d   
  via3  �d �x   
  via2  Yl Z   
  via2  f� Z   
  via2  ) �   
  via2  #�$ !   
  via2  K� #�x   
  via2  q� ��   
  via2  �� "�   
  via2  4, &
H   
  via2  � ��   
  via2  (!p �   
  via2  '�H o�   
  via2  ct 	�|   
  via2  &� ��   
  via2  � $�   
  via2  � ��   
  via2  
Zd ��   
  via3  Lp j�   
  via2  �� �   
  via2  ,p� �   
  via3  0� ��   
  via2  \� �   
  via2  iP n0   
  via2  <� @   
  via2  � j�   
  via2  �p ��   
  via3  �  �l   
  via2  &#� D   
  via2  �$ 	l   
  via2  )l 
f   
  via3  �4 ��   
  via2  g� $�   
  via2  "� %�(   
  via2  %`\ 	�T   
  via2  %ͼ �   
  via2  +8t �d   
  via3  *�l ��   
  via2  %� �h   
  via2  %
l �0   
  via2  �� �X   
  via2  d ��   
  via2  v� �   
  via2  &� ��   
  via3  � 9�   
  via3  � �   
  via2  �� !��   
  via2  	� �h   
  via2  *q< 	�|   
  via2  � n0   
  via2  �x �   
  via3  O\ �   
  via4  O\ �p   
  via4  � �p   
  via3  � �   
  via2  v( !QL   
  via2  �� $�H   
  via2  o �   
  via2  � 	Ѭ   
  via2  . D4   
  via2  ~< ��   
  via3  [ ��   
  via2  *�4 [<   
  via2  -�4 ��   
  via2  +� 	�T   
  via2  'g� �   
  via2  'o� ��   
  via3  GD 
 �   
  via2  | �l   
  via2  %�� �H   
  via   $�� �`   
  via2  #�� �X   
  via2  
�L ��   
  via2  � 9�   
  via3  d �   
  via2  =� gX   
  via2  � !*<   
  via2  � �   
  via3  d �   
  via3  d -   
  via2  %�| 	�,   
  via2  $y� 	�,   
  via   $y� 
�T   
  via2  3t �   
  via2  "P �   
  via2  '/@ C�   
  via2  '7 ��   
  via2  �� ��   
  via2  ;h "�    
  via2  �\ 	�\   
  via2  o ��   
  via2  0 �   
  via3  �� ��   
  via3  �� ��   
  via2  � ��   
  via2  �T 9�   
  via2  �d 
�D   
  via   *�t 4,   
  via2  )�$ �   
  via2  *<� 	E   
  via2  )�� �   
  via2  	�@ �   
  via2  4, ��   
  via3  d ��   
  via2  +֨ ��   
  via2  *�l �d   
  via2   @   
  via   �� �x   
  via    � �x   
  via2  ";� !�   
  via   !�  ʈ   
  via2  )_� �   
  via2   :  �   
  via2  -� �x   
  via3  ,4h ��   
  via3  ,4h �   
  via2  � #۰   
  via2  �D #۰   
  via2  �D $l8   
  via2  �� Al   
  via2  ` 9�   
  via3  ֌ 9�   
  via3  ֌ �   
  via2  	׈ !�   
  via2  �@ "�   
  via2  "� �x   
  via2  !?� �x   
  via   !?�  �   
  via2  $�, C�   
  via2  %;@ �   
  via2  �( `�   
  via2  �( 
B�   
  via2  `� k    
  via2  �$ ��   
  via2  �\ gX   
  via2  #z �   
  via2  �� �   
  via2  |� |   
  via2  �� "h�   
  via2  �� %    
  via2  \ T�   
  via2  _d �D   
  via2  << �D   
  via2  (�H    
  via2   6 �l   
  via3   �  �l   
  via3   �  h|   
  via2   �H h|   
  via    �H b|   
  via2  Ӝ �H   
  via2  :l ��   
  via   #  Sl   
  via2  � g�   
  via2  !	 ��   
  via2  !��  �l   
  via2   l�  �4   
  via2  	� #۰   
  via2  �\ !��   
  via3  E0 !��   
  via2  � %�(   
  via2  & ��   
  via2  �� ��   
  via   �l '   
  via   �\ '   
  via2  �d C�   
  via2  �� j�   
  via2  �� �X   
  via2  � �h   
  via2  �� ~�   
  via2  , C�   
  via2  � �   
  via2  �� ��   
  via2  �� ��   
  via2  �� �   
  via2  
� ��   
  via2  �� `�   
  via2  �� #۰   
  via2  �D !��   
  via2  b0 �   
  via3  �h !��   
  via3  �h !�8   
  via2  -	L j�   
  via2  ]L �   
  via2  �� �   
  via2  ��     
  via2  ^l ��   
  via2  � gX   
  via3  ]0 gX   
  via3  ]0 Ը   
  via2  �� !*<   
  via2  r� ��   
  via2  .M� j�   
  via3  -�� j�   
  via3  -�� ��   
  via2  "r\ �   
  via3  �� �   
  via3  �� �   
  via2   D %�8   
  via2  �� %�    
  via3  � %�    
  via2  	 � �    
  via2  � L�   
  via2   ��   
  via2  Q ��   
  via   Q ��   
  via2  � ��   
  via2  G  
�T   
  via2  �l $�   
  via2  p� !��   
  via2  #�� Al   
  via   "5� ��   
  via2  -4 �   
  via2  *ޜ [<   
  via   ,M� e    
  via3  ,�� ��   
  via4  ,�� ��   
  via4  -i  ��   
  via2  .L ��   
  via2  )�4 �p   
  via2  H�     
  via2  � o�   
  via2  !� |   
  via2  ^� ��   
  via2  W Y�   
  via3  ,� �   
  via2  #� �d   
  via2  � �x   
  via2  -*� ��   
  via2  �� %�   
  via2  �l �x   
  via2  �� 9�   
  via2  0 Al   
  via2  �H �   
  via2  + aX   
  via2  "f� &
H   
  via2   f� $݀   
  via2  �� 5�   
  via2  (�4 �0   
  via2  (� �@   
  via2  �� �d   
  via2  6d �   
  via2  �� ��   
  via   ., aX   
  via2  �8 Gh   
  via2   � k    
  via2  
� ��   
  via2  X� %�   
  via2  .� $�   
  via2  .� $%�   
  via3  .Y< $%�   
  via2  4� �x   
  via2   &�x   
  via2  -� ��   
  via3  ,� ��   
  via2  &o� ��   
  via2  $�L g�   
  via2   � �,   
  via2  �, j�   
  via2  ~ EP   
  via   zx e    
  via2  	�X  �   
  via2  � ��   
  via2  g� 8   
  via2  	Z� ʴ   
  via2  �L �D   
  via2  k� 	!�   
  via2  �p j�   
  via2  uL ��   
  via2  '� hx   
  via2  _� �l   
  via2  �� |   
  via2  D ��   
  via3  q� �d   
  via2  J� �d   
  via2  � !�8   
  via2  4 ��   
  via2  c0 �   
  via2  �� D0   
  via2  #�� Θ   
  via2  � 	E   
  via2  &X �p   
  via2  +� �x   
  via2  Z� �d   
  via2  �� 8   
  via2  	Z� !QL   
  via2  
, !�0   
  via2  &�� �    
  via2  �� �0   
  via2  � �   
  via2  *�� 8   
  via2  �H �   
  via2  T FL   
  via2  	A$ 9�   
  via2   �   
  via2  � ��   
  via2  �  �4   
  via2  �\ $�   
  via3  �\ !�8   
  via2  � T�   
  via2  2\ ��   
  via2  !�4 Al   
  via2   �� �|   
  via2  !l� @   
  via2  !I| �,   
  via2  0D Al   
  via2  4, ��   
  via2  � �x   
  via3  #� �8   
  via2  +�� 	u�   
  via2  
/l 8   
  via2  
7< �x   
  via2  %Ѥ 9�   
  via2  % �   
  via2  %� �   
  via3  )  �h   
  via2  @L `�   
  via2  � `�   
  via2  *@ #��   
  via2  *@ $l8   
  via2  �� %�8   
  via2  0� `�   
  via2  	� ��   
  via2  �d �   
  via2  `� dp   
  via2  �` ��   
  via2  ( 8   
  via   �� $   
  via2  +ax �x   
  via2  ʴ )�   
  via2  �< ��   
  via2  *�\ 9�   
  via   *�L 4,   
  via2  �  !�8   
  via2  � !�   
  via2  �� $�   
  via2  )<� sX   
  via2  *0� ��   
  via2  )� D   
  via2  S� �h   
  via2   � "p   
  via2  9P t�   
  via2  O� FL   
  via2  + D   
  via2  *y @   
  via2  K !tt   
  via2  Xl �0   
  via2  )�L k    
  via   |� �   
  via2  .� ��   
  via   ,*� e    
  via2  R$ �    
  via2  V �0   
  via3   �0   
  via3   )h   
  via2  8T &-p   
  via2  � &-p   
  via2  $jD �   
  via   #� <d   
  via2  P #��   
  via2  %J� %�(   
  via2  ~� ?�   
  via   [8 ��   
  via2  �  Gh   
  via2  #Q j�   
  via2  )� j�   
  via   *#    
  via2  H �x   
  via4  �, %�8   
  via2  �� 8   
  via2  +v� #��   
  via2  $�4 &   
  via2  q� �   
  via2  (� %�(   
  via2  6� D   
  via2  �L -   
  via2  /� ��   
  via2  � j�   
  via2  �\ Al   
  via2  }D 	�|   
  via2  �� Al   
  via   4� 	|   
  via2  $  !�(   
  via2  �0 #H   
  via2  }D o�   
  via   }D ��   
  via2  �� �   
  via2  ��     
  via4  %'� &�x   
  via2  %J� %��   
  via3  )�� ��   
  via2  *��  �\   
  via2  *�� ��   
  via2  *�� ��   
  via   *��    
  via2  Z�  �l   
  via2   X  �l   
  via2   X 2�   
  via3  
� %�8   
  via2  � "��   
  via2  �$ �0   
  via2  *�� �   
  via2  *�� ��   
  via2  &i� EP   
  via2  #� �8   
  via2  �� "��   
  via2  . !Md   
  via2  -O� �   
  via2  �t -   
  via3  |� -   
  via3  |� gX   
  via2  �� @   
  via2  l� �X   
  via2  �� �X   
  via2  �� �   
  via2  ƨ �X   
  via   ʐ �x   
  via2  *��  �l   
  via2  *p ��   
  via3  )�� ��   
  via2  � !�(   
  via2  �� !*<   
  via2   �, ��   
  via   U| '   
  via2   � ��   
  via2  -� \   
  via2  -�� K0   
  via3  -�� K0   
  via3  -�� 	p   
  via2  !h�  �\   
  via2  !`� ��   
  via2  *�� #$   
  via3  -�d D   
  via2  .&t D   
  via3  &� 9�   
  via2  �$ %�8   
  via2  Yl $�p   
  via3  |� $�p   
  via2  &�$ �   
  via2  &
H �4   
  via2  -�d D   
  via2  .� r@   
  via2  �� @   
  via   �x '   
  via2  �X �H   
  via   ۸ ��   
  via2  $�� :,   
  via2  $N� Θ   
  via3  $�� Θ   
  via3  $�� j�   
  via3  EP ��   
  via3  EP 	�,   
  via2  �4 �x   
  via2  �X !��   
  via3  �D !��   
  via3  �D #۰   
  via2  �4 �   
  via2  t� ��   
  via3  �� ��   
  via3  �� �   
  via2  Z� Al   
  via   �� b|   
  via2  1� �0   
  via2  ?� �x   
  via3  t �x   
  via2  �< ��   
  via2  � ��   
  via3  �� ��   
  via3  �� �h   
  via2  )P, ��   
  via2  !(H �   
  via3   �P �   
  via3   �P @H   
  via2  '� �   
  via2  M� ��   
  via2  � 2�   
  via2  E� 2�   
  via   E�    
  via2  &� o�   
  via2  r< ��   
  via2  + �h   
  via3  *� �h   
  via4  *� ��   
  via4  �� ��   
  via3  �� �h   
  via2  �� �x   
  via2  {, �h   
  via3  X �h   
  via2  $�\ @H   
  via2  .Y< ��   
  via3  .~X ��   
  via3  .~X ��   
  via2  
f %�8   
  via2  
m� %�    
  via3  
� %�    
  via2  �� �l   
  via2  �P �   
  via2  ׄ �   
  via2  EP k    
  via3  &�D �   
  via3  '}`  ��   
  via4  '}`  ��   
  via4  )�0  ��   
  via3  )�0 |   
  via2  %�<  �\   
  via2  �� 2�   
  via2  0� �   
  via2  - @   
  via2  %�� 	�T   
  via2  #�� ��   
  via4  #G@ $�   
  via4  $�D $�   
  via3  $�D #۰   
  via2  &; ��   
  via2  �� �   
  via2  "d� j�   
  via2  �X ��   
  via2  ')d el   
  via2  < |   
  via2  |l ��   
  via2  	0 ��   
  via2  .?� #۰   
  via3  -�� #۰   
  via4  -�� $�   
  via4  .6 $�   
  via4  � ��   
  via3  �\ $�   
  via2  �H #��   
  via2  r� �x   
  via4   @ �x   
  via3   @ �h   
  via2  �4 �h   
  via2  &�� BD   
  via2  '�t ��   
  via2  r� $�   
  via3  N ��   
  via2  �� �   
  via2  +d !�8   
  via2  #� #۰   
  via3  #G@ #۰   
  via2  � !�8   
  via2  QP �x   
  via2  4p ��   
  via2  '\, 	!�   
  via4  $�L '�   
  via2  (� #��   
  via2  �,  �   
  via2  � �   
  via3  9 �   
  via4  9 ��   
  via4  � ��   
  via3  � �   
  via2  *d !�(   
  via2  '� !��   
  via2  Μ    
  via3  +�\ `�   
  via4  +�\ �L   
  via4  )�� �L   
  via2  +� ��   
  via4  v� �h   
  via3  v� �x   
  via2  �     
  via2  !,     
  via2  !, k    
  via2  �� �   
  via2  �t 	�,   
  via3  � 	�,   
  via4  � 	    
  via4  j� 	    
  via2  SD �   
  via2  +\ !�8   
  via2  I� 8   
  via2  + �   
  via2  .*\ ��   
  via2  *� �   
  via2  K 2�   
  via2  	�  ,�   
  via3  	'�  ,�   
  via4  	'�  S�   
  via4  ��  S�   
  via3  ��  ,�   
  via   O� ��   
  via2  �D :,   
  via2  (�� �   
  via2  +�$ `�   
  via3  �� ��   
  via4  �� ��   
  via4  �� ��   
  via2  )V 	�,   
  via2  $�� 	!�   
  via2   @ 	l   
  via2  �8 �   
  via2  m� &
H   
  via2  �� -   
  via2  �D |   
  via2  )@� Ml   
  via2  : �    
  via2  � !�   
  via2  #� !�(   
  via2  +\ !�(   
  via2  � ��   
  via2  &�� \   
  via2  #� 	�T   
  via2  �l �h   
  via2  Y� �d   
  via2  �, |   
  via2  "Ep f   
  via2  �0 %�(   
  via2  *mT Y$   
  via2  � `�   
  via2  &�, k    
  via2  %q� �   
  via3  '�� �   
  via2  �  �   
  via2  l� ��   
  via2  j� �   
  via2  �\ %�    
  via2  ;� #۰   
  via2  '0 	l   
  via2  '� 	h4   
  via2  '� 	�,   
  via2  �\ &
H   
  via2  �D %�8   
  via2  [� %�8   
  via2  [� %�    
  via2  e�    
  via2  � ��   
  via3  b0 ��   
  via3  b0 ��   
  via2  �d Al   
  via2  g� !��   
  via2  N ��   
  via2  %'� ��   
  via2  �l ��   
  via2  S� �X   
  via2  bx %�8   
  via2  bx &
H   
  via2  $�D ��   
  via2  &` L�   
  via2  �� &
H   
  via   �p 0D   
  via2  q� 	�,   
  via2  ,�� �    
  via2  �� ��   
  via2  )H ��   
  via3  ˈ �X   
  via2  �� \   
  via2  
90 �   
  via2  
= -   
  via2  	�� Al   
  via2  � h|   
  via2  zx �0   
  via2  zx @   
  via2   �   
  via2  LH j�   
  via2  v$ 9�   
  via2  �H �   
  via2   �  �l   
  via2  �  �\   
  via2  D� !�(   
  via3  -&� `�   
  via2  �� !��   
  via2   � j�   
  via3  �� ۔   
  via2  � 
F�   
  via2  �� \   
  via2  )�D ��   
  via2  �l ��   
  via2  *H8 \   
  via2  	P� o�   
  via3  &� 4   
  via2  �l "`   
  via2  �� Ј   
  via2  %� D   
  via2  %x u   
  via2   4 ��   
  via2  m\ o�   
  via2  u, !�8   
  via2  �L %�8   
  via2  	T� $�   
  via2  !	 #$   
  via2  �� !�8   
  via2  &Z\ �0   
  via2  �  &-p   
  via2  �� ��   
  via2   \ 	�,   
  via2  "�� #�x   
  via2  r� $�   
  via2  _� D   
  via2  � k    
  via2  %'� %��   
  via3  $ی %��   
  via4  $ی &�x   
  via2  *<� |   
  via2  $�4 'F�   
  via3  $�\ 'F�   
  via4  $�\ '�   
  via2  �d $�   
  via2  �X !�8   
  via2  "9� 9�   
  via2  �l �   
  via2  �� #$   
  via2  +cl `�   
  via2  �0 ��   
  via2  �  4   
  via4  #t, &�x   
  via2  �� ��   
  via2  _$ 9�   
  via2  o  ,�   
  via3  ��  ,�   
  via4  ��  S�   
  via4  ��  S�   
  via3  �� |   
  via2  x 	l   
  via2  ` 	�T   
  via2  �X ��   
  via2  #I4 %��   
  via3  #l\ %��   
  via4  #l\ &^D   
  via2  +� #۰   
  via2  :� `�   
  via2  {L `�   
  via2  hx |   
  via3  W Y�   
  via2  K� k    
  via2  �� �X   
  via2  �, j�   
  via2  =� k    
  via2  �� �   
  via2  �� ��   
  via2  l� k    
  via2  *6� �h   
  via2  (�� 8   
  via2  v� :,   
  via2  p� ��   
  via2  (�$ Al   
  via2  "`� �   
  via2  �p �   
  via2  	�L #$   
  via2  �� �X   
  via2  #�� ��   
  via2  �� `�   
  via2  w� !�8   
  via2  (
  EP   
  via2  'k� -   
  via2  �� �x   
  via2  0� Ј   
  via2  k� "�   
  via2  @� jp   
  via2  �� �h   
  via2  \ @   
  via2  � j�   
  via2  �P h|   
  via3  �p h|   
  via3  �p 5�   
  via2  ؀     
  via2  "��     
  via2  %� 	l   
  via   8 ��   
  via2  �h D   
  via2  LL ��   
  via2  �� �x   
  via2  R� \   
  via2  R� Al   
  via2  � �4   
  via2  	� �   
  via2  ,m ��   
  via2  +�P �x   
  via2  L |   
  via2  n4  �\   
  via2  �, |   
  via2  �� n0   
  via2  )0� 	�T   
  via2  !&T D   
  via2  !,0     
  via2  �t aX   
  via2  �@ Ј   
  via2  ,v� �h   
  via2  ,v� �X   
  via2  ø �   
  via2  �� #$   
  via2  a D4   
  via2  �L ��   
  via2  ��    
  via3  :� =`   
  via2  �    
  via   �  0D   
  via2  H |   
  via2  'H� 9�   
  via2  �\ 5�   
  via2  &�  ��   
  via2  (T8 BD   
  via2  "?� %�@   
  via2  !� $�   
  via2  �t T�   
  via2  $ � �   
  via2  %�� �   
  via2  "7� ��   
  via2  -�     
  via2  ,M� ��   
  via2  2� �   
  via2  "� ��   
  via   � aX   
  via2  �  &
H   
  via2  ��    
  via2  �0 !�8   
  via   �� 
�,   
  via2  	�t ��   
  via2  �� �   
  via2  � #$   
  via2  +�P k    
  via2  i� �   
  via2  m� P0   
  via2  )8� �X   
  via2  "9� Al   
  via2  �$ 	l   
  via2  �� ��   
  via2  $� ��   
  via2  � ��   
  via3  6� ��   
  via3  ڼ 	l   
  via2  5� C�   
  via2  =� j�   
  via2  )�4  �l   
  via2  *4 ��   
  via2   WL 
ϔ   
  via2  #�� 	�,   
  via2  '�4 $�   
  via2  )R  #۰   
  via2  �0 ��   
  via2  � 	l   
  via3  y 	l   
  via3  y 	�,   
  via3  '�4 n�   
  via2  &�, �\   
  via2  $
� �   
  via2  $
� -   
  via3  �� ��   
  via2  ;D $�   
  via2  +�P D   
  via2  �X �d   
  via2  #�` 	E   
  via2  �$ %�8   
  via2  �� &-p   
  via   � �x   
  via2  +Դ ��   
  via2  #��    
  via2  S� #$   
  via2  �� ��   
  via2  � ""H   
  via2  &� %�    
  via2  +,� ��   
  via2  #Q D   
  via2  
m� o�   
  via2  �� ��   
  via2  (�� p�   
  via2  -�d L�   
  via2  �L �X   
  via2  �� 	E   
  via2  &�\  ��   
  via2  �� ��   
  via2  %C 4   
  via4  &�  ��   
  via4  &�D  ��   
  via2  �4 ��   
  via2  �X ��   
  via2  �� j�   
  via2  � �x   
  via2  � D   
  via2  �X ��   
  via2    �\   
  via2  �� k�   
  via4  6� 	!�   
  via2  �l ɔ   
  via2  � ��   
  via2  %H P0   
  via2  'Z8    
  via2  \ %�8   
  via2  x@ &
H   
  via3  Lp ��   
  via2  y\ ��   
  via2  ,Ҝ �x   
  via2  �, �   
  via3  !� ��   
  via2  '� p�   
  via2  	�T 	!�   
  via3  Kt 	��   
  via2  �� \   
  via3  @L `�   
  via2  zT �4   
  via4  $;d �(   
  via2  %�� @   
  via2  �� <�   
  via2  � ��   
  via2  ,�$ -   
  via2  �� )h   
  via2  P ��   
  via2  �� �   
  via2  -0  �l   
  via2    �l   
  via3  �� gX   
  via3  �� @H   
  via2  -"� j�   
  via2  �� k    
  via2  
�, ��   
  via   .X R�   
  via2  ,*� ��   
  via3  �$ �X   
  via2  !� o�   
  via3   �` �D   
  via2  #ݤ ��   
  via2  4 �h   
  via2  2 j�   
  via2  	�� 	�,   
  via2  �� Al   
  via2  �� �h   
  via2  )�  ��   
  via2  ";� �X   
  via2  $� !�   
  via2  , &
H   
  via2  1� &
H   
  via2  �\ !�   
  via2  {p @H   
  via2  X 8   
  via2  _@ ��   
  via2  | ��   
  via2  *# ��   
  via2  (m� j�   
  via2  � !�8   
  via2  �l gX   
  via2  �� -   
  via2  �� ��   
  via2  �� �h   
  via2  $T �h   
  via2  )�� �h   
  via2  )  @   
  via2  �� %�8   
  via2  � %�(   
  via3  )X �   
  via2  $� ��   
  via2  (B� �h   
  via2  '�� �X   
  via2  :L #۰   
  via2  "�8 !�8   
  via2  k� !f�   
  via2  ��  �4   
  via2  �  �\   
  via2  �  �\   
  via2  3�  �\   
  via2  D ��   
  via2  N �x   
  via2  �l     
  via2  �� C�   
  via2   	l   
  via2  �X ��   
  via2  $�$  �l   
  via2  $H  �\   
  via2  $�$ �0   
  via2  $�X �x   
  via3  ^H A�   
  via2  ژ #$   
  via2  � ��   
  via2  �� `�   
  via2  �� �   
  via2  �X  �\   
  via2  �D �|   
  via2  VX �   
  via2  � �   
  via2  � ��   
  via2  @H L�   
  via2  '� o�   
  via2  ""H 	�,   
  via2  �X 	E   
  via2  ] �D   
  via2  � �   
  via2  %/� �   
  via2  �� @   
  via2  ,�< &
H   
  via2  �� o�   
  via3  Y� ��   
  via2  /  j�   
  via2  #�� �   
  via2  !`� �   
  via2  �L  �\   
  via2  :� ��   
  via2  '� 	�T   
  via2  
� \   
  via2  	�� \   
  via2  � \   
  via2  P4 D   
  via2  ~� D   
  via2  4L C�   
  via2  �p Al   
  via2  ��     
  via2  .�L -   
  via2  �� �   
  via2  O8 �   
  via2  )�L -   
  via2  '\, >0   
  via2  % Ј   
  via3  %A Ј   
  via4  %A e@   
  via4  &�� e@   
  via2  (�� �h   
  via2   f� !�   
  via2  !� ��   
  via2  !� `�   
  via   �� 
�,   
  via2  � h|   
  via2  � ��   
  via2  �� 	�T   
  via2  +�� Al   
  via2  +Դ h|   
  via2  -�` 	p   
  via2  ,�L D   
  via2  � �h   
  via2  �� @   
  via2  L $��   
  via2  @L $�   
  via2  &�, #��   
  via2  &Ǽ !�   
  via2  �l f�   
  via2  �� @   
  via2  )� 	l   
  via2  )�l 	�,   
  via2  qd ��   
  via2  �� ��   
  via3  &-p 
#�   
  via2  #EL :,   
  via2  W !�   
  via2  �  #��   
  via2  �H C�   
  via2  �0 j�   
  via2  �p !�(   
  via2  	�p @H   
  via2  �� ��   
  via2  �D ��   
  via2  �� k    
  via2  I� k    
  via2  (+4 �p   
  via2  #x `�   
  via2  )  ��   
  via2  &� ��   
  via3  &ό ��   
  via4  &ό �   
  via4  '�l �   
  via2  �� j�   
  via2   E�  �l   
  via2  *�8 �   
  via2  *�8 ��   
  via2  �<  �\   
  via2  _  o�   
  via2  $  #$   
  via2  $�� �H   
  via2  .6 �   
  via2  � #$   
  via2  �� ��   
  via2  "\� 9�   
  via2  %ͼ C�   
  via   +�� b|   
  via2  *u$ ��   
  via2  "�d @   
  via2  +d �h   
  via2   6 ��   
  via2  4l    
  via2  $�( �x   
  via2  $� �h   
  via2  ,<8 �   
  via2  �x ��   
  via2  \ 	E   
  via    b|   
  via2  �4 h|   
  via2  ְ 	l   
  via2  �\ 	�,   
  via2  ݄ �   
  via2  9t h|   
  via2  cP #��   
  via2  � !�(   
  via2  <� ��   
  via2  
�X ��   
  via2  )�� @H   
  via2  (�� ��   
  via2  %� k    
  via3  � �   
  via2  �, |   
  via2  �� !�(   
  via2  0� !�8   
  via2  �� gX   
  via2  3t !�8   
  via2  '�� @H   
  via2  %w� gX   
  via3  &X �p   
  via2  28 	E   
  via2  � ��   
  via2  �t ��   
  via2  �0 @H   
  via2  � &
H   
  via2  'k� �h   
  via2  *2� �    
  via2  �� ��   
  via2  �  ��   
  via2  �T �   
  via2  �H `�   
  via2  
� k    
  via2  �� �   
  via2  Yd �   
  via2  �� ��   
  via2  �� �   
  via2  �� �   
  via2  )mx @H   
  via3  �4 	�,   
  via2  T� ��   
  via2  I ��   
  via2  .;� �x   
  via2  -[T @H   
  via2  D gX   
  via2  ܬ -   
  via2  �� �   
  via2  ,aT !�(   
  via2  �� �    
  via2   Ȕ �x   
  via2  ,]l 8   
  via2  �T �   
  via2   � Ј   
  via2  !� �   
  via2  �� 	�,   
  via3  J0 	�,   
  via4  J0 ��   
  via4  �4 ��   
  via2  �  �l   
  via   � $   
  via2  � D   
  via2  y 	�,   
  via2  �� !�   
  via   �   @   
  via2  �x !�   
  via2  "� �x   
  via2  ܌ Ј   
  via2  *D 	l   
  via3  �4 	l   
  via2  W0 j�   
  via2  �\     
  via2  ۸ 	l   
  via2   \ 	E   
  via2  "�� �   
  via2  )	� 	E   
  via2  ! j�   
  via2  � ��   
  via2  )<� !�8   
  via2  
�� H�   
  via2  Nd �x   
  via2  l� Al   
  via2  �X ��   
  via2  ;l C�   
  via2  c� Al   
  via2  [X ��   
  via2  &; h|   
  via2  &; Al   
  via2  (�� .,   
  via2  *�L Al   
  via2  !A� #��   
  via2  !�� %�(   
  via2  ,t� :p   
  via2  ,� D   
  via2  , �0   
  via2  , @   
  via2  �� P   
  via2  	-� @   
  via2  �� %    
  via2  � &
H   
  via2   8   
  via2  �0 @H   
  via2  � 8   
  via2  N� �0   
  via2  	bX !�8   
  via2  �� �   
  via2  �� -   
  via2  �� #۰   
  via2  �� $�   
  via2  � %�(   
  via2  'b ��   
  via2  Ml !�   
  via2   #��   
  via2  #nP 	l   
  via2   6 ��   
  via3  *0� ��   
  via2  '�� !�   
  via2  � 6�   
  via2  	��  �\   
  via2  (�� ��   
  via2  (Ì ��   
  via2  
\ �    
  via2  	bX ��   
  via2  "?� #۰   
  via2   � #��   
  via2  � %�8   
  via2  !� &
H   
  via2  � v    
  via2  x j�   
  via2  0 @H   
  via2  a4 j�   
  via2  , ��   
  via3  \�  �\   
  via2  XL |   
  via2  �� 	�T   
  via2  e  	E   
  via2  
? &
H   
  via2  �  �l   
  via2  (3 �   
  via2   � ��   
  via2  	� l   
  via2  �X ��   
  via2  ' 	E   
  via2  � �0   
  via2  ��     
  via2  T� �h   
  via4  Yl �,   
  via2  |L #$   
  via2  #� �h   
  via2  �� �h   
  via2  }� �X   
  via2  �� 8   
  via3  �< �0   
  via2  -, �    
  via2  �4 �x   
  via2  �, �h   
  via2  ,�� !�   
  via2  ?t �H   
  via2  $� -   
  via2  $^� �    
  via2  
�� |�   
  via2  h� �   
  via2  4� #۰   
  via3  (�� �@   
  via2  (B� @H   
  via2  Q ��   
  via2  "�x %�8   
  via2  �� %�(   
  via2  �l     
  via2  
3T D   
  via2  AH �(   
  via2  �� ��   
  via2  ��     
  via4  
  ��   
  via2  �� ��   
  via2  !� ��   
  via2  +iH o�   
  via2  *�� @   
  via2  �� 9�   
  via2  �� `�   
  via2  D4 	�,   
  via2  �� 	�,   
  via2  �d #$   
  via2  y\ �   
  via2  7 �    
  via2  �$ ��   
  via2  	�� ��   
  via2  9� �X   
  via2  �� ��   
  via2  �\ C�   
  via2  � �   
  via2   D �0   
  via2  �H %�(   
  via2  �H ��   
  via2  � 	E   
  via2  6� 	l   
  via2  � ��   
  via2  B� Al   
  via2    ��   
  via2  �D 9�   
  via2  
;$ C�   
  via2   ;� ��   
  via2  o  �l   
  via2  y� �h   
  via2  � j�   
  via   $ � 
�,   
  via2  �� C�   
  via2  +X 8   
  via2  (4�  �\   
  via2  �� ��   
  via2  �  �\   
  via2  Y$ h|   
  via2  �� \   
  via2  � �T   
  via2  �` �   
  via2  -� �|   
  via2  '�� .,   
  via2  "� C�   
  via2  � j�   
  via2  D ��   
  via2  	�� "��   
  via2  � !�   
  via2  #1� g8   
  via2  θ ��   
  via2  �� D   
  via2  #� ��   
  via2  .�� �0   
  via2  -E� j�   
  via2  :, �   
  via2  +B8 8   
  via2  -j� ��   
  via2  !� ��   
  via2  $�� ��   
  via2  (�� ��   
  via2   d� \   
  via2  -�� 8   
  via2  +�L @H   
  via2  +�� ��   
  via2  +�� j�   
  via2  !� 
j   
  via2   � Al   
  via2  *� �   
  via2  4� �    
  via2  �� h|   
  via2  C� o�   
  via2  �� ]T   
  via2  :� |   
  via2  � `�   
  via2  8 ��   
  via2  � @H   
  via2  :l gX   
  via2  �t 8   
  via2  &�� gX   
  via2  &� 8   
  via2  �0 !�   
  via2  � �x   
  via2  #� #H   
  via2  +�4 !�   
  via2  -�t !�(   
  via2  #I4 �    
  via2  Ƥ �    
  via2   >   
  via2  D j�   
  via2  @$ ��   
  via2  _� �X   
  via2  	Ք ��   
  via2  ;� ��   
  via2  �� �D   
  via2  �4 ��   
  via2  �T 9�   
  via2  �4 T�   
  via2  �� ��   
  via2  � ��   
  via2  %�D  �l   
  via2  !�d �0   
  via2  �t j�   
  via2  o �h   
  via2  ?t �h   
  via2  �  _@   
  via2  4 �h   
  via2  �l #��   
  via2  &�� ��   
  via2  &��    
  via2  � Ј   
  via2  �, $�   
  via3  '�l ��   
  via2  (�� ��   
  via2  (Jt ��   
  via2  &�� j�   
  via2  � !�(   
  via2  � !�   
  via2  � |�   
  via2  k�  �\   
  via2  � |�   
  via2  ct |   
  via2  $f\ �h   
  via2  g\ ��   
  via2  U� Al   
  via2  Rp @H   
  via2  
�l j�   
  via3  *� )h   
  via2  '�l o�   
  via2  -g �x   
  via2  U� gX   
  via2  [� aX   
  via2  � gX   
  via2  +�D �   
  via2  ܈ $�   
  via2  Xl %�(   
  via2  |L �   
  via2  "� �h   
  via2  k #��   
  via2  �� #��   
  via2  �d #۰   
  via2  �\ 0�   
  via2  � %�(   
  via2  i �   
  via2  S$ #۰   
  via2  �  ��   
  via2  &R� ��   
  via   �� ��   
  via2  &N� ��   
  via2  K� !�(   
  via2  � #��   
  via2  (a� j�   
  via2  +�� 	l   
  via2  %s� �0   
  via2  %� 8   
  via2  6� @H   
  via2  d$ @H   
  via3   �( �p   
  via2  +�L �h   
  via2  �| ��   
  via2  L !�   
  via2  � gX   
  via2  � @H   
  via2  &q� @H   
  via2  �� @H   
  via3  -�� ��   
  via2  +s �   
  via2  �� |�   
  via2  ֬     
  via2  �� %�8   
  via2  � %�8   
  via2  "�l    
  via2  �P &P�   
  via2  � #۰   
  via2  � ��   
  via2  �0  �l   
  via2  r� ��   
  via2  '� o�   
  via2  �� %�8   
  via2  r� %�(   
  via2  d %�8   
  via2  �� j�   
  via2  
�� C�   
  via3  L |   
  via2  `�  �\   
  via2  
�| T�   
  via3  -j� ��   
  via2  +�� h|   
  via2  %)� h|   
  via2  
-x �h   
  via2  	)� �   
  via3  �, d�   
  via2  �,    
  via4   | <   
  via2  �, `�   
  via2  �< &-p   
  via2  x� ��   
  via2   �� �   
  via2  O� �x   
  via2  )� �x   
  via2  '�l ��   
  via2  �� &
H   
  via2  �� #۰   
  via2  (RD �x   
  via2  (V, Ј   
  via2  ' ��   
  via2  #�� �x   
  via2  ! �   
  via2  l �    
  via2   �d f   
  via2  �� �   
  via3  XL |   
  via2  %� @H   
  via2  ,�� Al   
  via2  �l ��   
  via2  -v� k    
  via2  �� f   
  via2  (� �   
  via2  kD �x   
  via   +:h  ʈ   
  via2  �� #۰   
  via2  �� ��   
  via2  H� %�(   
  via2  "Gd ��   
  via2   �� ��   
  via2  !� �h   
  via2  ";� 8   
  via2  �  �   
  via2  Ŭ  �\   
  via   � ��   
  via2  �, j�   
  via2  �0 �   
  via2  �� �   
  via2  � 9�   
  via2  (, �   
  via2  � Al   
  via2  x� \   
  via2  - d   
  via2  ׬ �   
  via2  $u� !�8   
  via2  , o�   
  via2  *S� �    
  via2  &$ �h   
  via2  #b� �h   
  via2  Ј ��   
  via2  c� ��   
  via2  �$ ��   
  via2   
ϔ   
  via2  ��  �l   
  via2  �� |   
  via2    8   
  via2  +�p    
  via2  �l "��   
  via2  l� �0   
  via2  
� !�0   
  via2  \0 �   
  via2  t j�   
  via2  $�X 8   
  via2  |� ��   
  via2   �h   
  via   !�  �   
  via2  ;� �0   
  via2  �\ #۰   
  via2  gX #��   
  via2   .H k    
  via2  �p �   
  via2  � !�(   
  via2  !� @H   
  via2  v %�@   
  via2  
�� %�8   
  via2  � $L�   
  via2  �� "��   
  via2  !�� $�   
  via2  �� ��   
  via3  �P #$   
  via2  �� 	�\   
  via2  	P� �0   
  via2  	� �    
  via2  � "�    
  via2  �0 %�8   
  via   �� ��   
  via2  �p D   
  via2  %A 	E   
  via2  X �h   
  via2   � @   
  via2  (�� 	l   
  via2  &� ��   
  via2  7� #۰   
  via2   � ��   
  via2  
�x 	l   
  via2  V4 	E   
  via2  SD Al   
  via2  �� ��   
  via2  �x 	l   
  via2  c, !�    
  via2  $ #۰   
  via2  H� ��   
  via2  � %�(   
  via2  Ԙ "(   
  via2  $ ��   
  via2  !Md Θ   
  via2  �  	l   
  via2  � 	E   
  via2  1 	l   
  via2  #5�  �\   
  via2  -A� �   
  via2  +�< -   
  via2  Z<    
  via2  s| ��   
  via2  � �   
  via2  �� ��   
  via2  �< -   
  via2  ȼ �    
  via2  �$ �0   
  via2  � �x   
  via2  � %�8   
  via2  �� ��   
  via2  Ԙ j�   
  via3  &�� >0   
  via2  &o� !�(   
  via2  !l� �,   
  via2   �� ��   
  via2  �` ��   
  via2  Ќ o�   
  via2  7� 8   
  via2  �� |   
  via2  �� 	�d   
  via2  !
� C�   
  via2  �L ��   
  via2  >T ��   
  via2  %�H !�   
  via2  (>� !�8   
  via2  �� @H   
  via2  (L �X   
  via2  +e` !�(   
  via3  � ��   
  via2  � �0   
  via   �  '   
  via2  /  �h   
  via2  �T $�   
  via2  #�  C�   
  via3  $� �x   
  via2   C� �0   
  via2  ,�D o�   
  via2  Mh $�`   
  via2  
�h �   
  via2  �� �h   
  via4  P� w@   
  via2  � �x   
  via2  �@ ""H   
  via2  �� �0   
  via3  ,0� �   
  via2  #` �0   
  via2   j� @H   
  via2  �` �x   
  via   #�� <d   
  via2  %'� D   
  via2  � �X   
  via2  � ��   
  via2  *�d P0   
  via2  &�� @H   
  via2  ,�< �h   
  via2  Lp ��   
  via2  �� j�   
  via2  �� `�   
  via2  �T 9�   
  via2  (�  �l   
  via2  $�D  �l   
  via2  �� D   
  via2  *P �X   
  via2  (�� �h   
  via3  (]� �    
  via2  *�� 	l   
  via2  " :,   
  via2  
� ��   
  via2  )�X L�   
  via2  6�  �\   
  via2  k$ ��   
  via2  (t  �l   
  via2  �  �   
  via2  ô U`   
  via2  � x�   
  via2  L 	l   
  via2   ��   
  via2  	� ��   
  via2  
 � ��   
  via2  /$ ׬   
  via2  	w� o�   
  via2  �� �0   
  via2  � �h   
  via2  %�$ $%�   
  via2  !E� #۰   
  via2  �� j�   
  via2  a� ��   
  via2  x� $'�   
  via2  � %�(   
  via2  �� Ј   
  via2  � %�(   
  via2  l�  ��   
  via2  � !�8   
  via2  � 9�   
  via2  d �,   
  via2  d �,   
  via2  e$ 9�   
  via3  8 n�   
  via2  
�� ��   
  via2  ~d �   
  via3   a @H   
  via2  +܄ �x   
  via2  �D #۰   
  via2  6� #��   
  via2  "�� �x   
  via2  �t ��   
  via2  Y$ �   
  via2  '0  �l   
  via2  5$  �l   
  via3  0� dH   
  via2  %Ѥ \   
  via2  ,0� ��   
  via2  +�� �    
  via3  ,p� �`   
  via2  ,*�     
  via2  ! %�8   
  via2  ( ��   
  via2  � `�   
  via3   "��   
  via2  >� #۰   
  via3  g� &�x   
  via2  #D %�8   
  via4  � !�8   
  via2  N� !�(   
  via2  �T !�(   
  via2  R �x   
  via3  ,Ҝ Ը   
  via2  #�D @H   
  via2  !�L ��   
  via2  �� �   
  via2  e  !�   
  via3  2� ��   
  via2  � �   
  via3  *�l �d   
  via2  �� @   
  via2  � &
H   
  via3   ;� �   
  via2  (c� Ml   
  via2  .d� Al   
  via2  )'( Al   
  via2  '� �   
  via2  ,δ \   
  via2  
p  �l   
  via2  � Al   
  via2  ܰ 9�   
  via2  
� �X   
  via2  @l $��   
  via2  � !�   
  via3  +�� @   
  via2  +(� �0   
  via2  � ��   
  via2  �\ h|   
  via2  �L @H   
  via2  r@ gX   
  via2  Al &-p   
  via2  &\ &
H   
  via2  �$ �h   
  via2  %8 j�   
  via2  �� �0   
  via2  
�� #۰   
  via2  Ь ��   
  via2  Ԙ !�(   
  via2  )�� !��   
  via2   �P %�(   
  via2   ��   
  via2  5�  �\   
  via2  �� Al   
  via2  g\ =`   
  via2  3 	l   
  via3  $  #$   
  via2  '�, ��   
  via4  "�  �   
  via2  # 0 �   
  via2  !� %�8   
  via2  'k� ��   
  via2  � D   
  via2  � @H   
  via2  N� ��   
  via2  �� \   
  via2  -,  �\   
  via2  +S� 	�,   
  via2  %� �h   
  via2  
� P   
  via2  ( j�   
  via3  Yl Z   
  via2  %�4 ��   
  via2  _d sX   
  via2  � �   
  via2  �� Ј   
  via2  �� 8   
  via2  p 9�   
  via   "� b|   
  via2  ְ  �l   
  via2   :,   
  via2   �   
  via2  @ 	Ѭ   
  via2  �P #$   
  via2  �� ��   
  via2  �L  �\   
  via2  )� ��   
  via   W� 	|   
  via2  	�� ��   
  via2  
�l  �\   
  via2  �� |   
  via2  _$ �H   
  via2  *�d �x   
  via2  o !�(   
  via2  '�� ��   
  via2  %dD �x   
  via2  L� 
B�   
  via2  Q� Al   
  via3  (�$ -   
  via2  ]p 	E   
  via2  �4 !�8   
  via2  '��     
  via2  &h �   
  via2  )�0  �\   
  via2  n� |   
  via2  >� j�   
  via2  ?P #۰   
  via2  -ȴ D   
  via2  ,ք 	l   
  via   ."� ��   
  via2  , Al   
  via2  �� !�8   
  via2  � �0   
  via2  -Wl  �   
  via2  )� �   
  via2  �� �   
  via2  �x �   
  via2  $�� 9�   
  via2  L ��   
  via2  � D   
  via3  � `�   
  via2  (@� ��   
  via2  , 9�   
  via2  �� �   
  via2  �� ��   
  via2  �� 
(   
  via2  � �   
  via2  qd �`   
  via2  
'� ��   
  via2  '-L "A�   
  via2  #EL !�(   
  via2  1� f�   
  via2  q� ��   
  via2  _� �   
  via2  \0 Al   
  via2  #�4  �l   
  via2  '�L  �l   
  via2  *W� D   
  via2  "�, �   
  via2  $=X ��   
  via2  > %�(   
  via2   ;� %�8   
  via2  "�4 �   
  via2  (D� �   
  via2  '-L u   
  via2   UX D   
  via2  �H 	��   
  via2  U` 	l   
  via2  
�� |   
  via2  � ��   
  via2  � �    
  via2  � C�   
  via2   h|   
  via2  K� ��   
  via2  	� ��   
  via2  �� ��   
  via2  	� ��   
  via2    �\   
  via2  � �x   
  via2  �� j�   
  via3  #D %�8   
  via2  �X !�(   
  via2  )�| ��   
  via2  -e �   
  via4  N� !Ĉ   
  via2  �� @H   
  via   H  ʈ   
  via2  V0 D   
  via2  ô     
  via2  �� �   
  via2  	h4 8   
  via2  ̤ P0   
  via2  z4 ��   
  via2  � $%�   
  via2  !tt !�   
  via2  � !�(   
  via3  'T ��   
  via2  &�� >0   
  via2  #�� �x   
  via2  $� �x   
  via2   � !��   
  via2  �� !�   
  via2  &Vt o�   
  via2  $�X "��   
  via2  $C4 #��   
  via2  %
l #��   
  via2  &� #��   
  via2  � o   
  via2  4     
  via2  �� j�   
  via2  t4 C�   
  via2  $  %�   
  via2  /� j�   
  via2  x j�   
  via2  ct C�   
  via2  !Md ��   
  via2  "nt  �\   
  via2  . ��   
  via2  +M� 9�   
  via2  ){$ 	A$   
  via2  +u  �   
  via2  *�d �D   
  via2  #;� ��   
  via2  k� l   
  via2  !x �h   
  via2  �L Y�   
  via2  �x �   
  via3  X �x   
  via2  � @H   
  via   (� �x   
  via2  �� �0   
  via2  '�d ��   
  via2  �8 5�   
  via2  e� &-p   
  via2  Ը �h   
  via2  	��  	�   
  via2  ��  �\   
  via2   � !�(   
  via2  �  o�   
  via2  "�d !�   
  via2  $�� !�   
  via2  &�� )h   
  via2   G� #$   
  via3  )�  ��   
  via2  )�� �X   
  via2  U� ��   
  via2  �� ��   
  via2  �� 2�   
  via2  -0 ��   
  via2  $G �   
  via2  )� 9�   
  via3  +	� -   
  via2  *�� �   
  via2  �< #$   
  via2  t �   
  via2  �  �\   
  via2  �  �l   
  via2  ' P0   
  via2  |� !�   
  via2  !p� k    
  via2  �8 	l   
  via2  �� ,   
  via2  #d� #$   
  via3  .*\ ��   
  via2  )g� ��   
  via2  %�� �   
  via2  w �   
  via3  �, m�   
  via2  +�� ��   
  via2  -�H L�   
  via2  -G� ��   
  via2   4$ ��   
  via2  %� ��   
  via2  + �   
  via2  (�� k    
  via2  l� 	�,   
  via2  7� 9�   
  via2  ($  S�   
  via2   �� ��   
  via2  "� !�(   
  via2  x� @H   
  via2  �, "�   
  via2  E0 #۰   
  via3  '!� j    
  via2  &1X �    
  via2  %�d ��   
  via2  '�p j�   
  via2  (� o�   
  via2  ( �h   
  via3  'VP f   
  via2  *a� �   
  via2  )�d ��   
  via2  K0 @H   
  via3  t �0   
  via2  �p �    
  via2  �X �x   
  via2  =� !�(   
  via2  �4 \   
  via2  �0 9�   
  via2  ˈ `�   
  via2  �� 9�   
  via2  � 
�l   
  via2  �0 ��   
  via2  �H ��   
  via2  ,X �X   
  via2  :L ��   
  via2  �p �0   
  via2  � !*<   
  via2  D �   
  via   ��  ʈ   
  via2  � ��   
  via2  �� 8   
  via2  4 �h   
  via2  �� >   
  via2  /D �   
  via2  *# �   
  via2  "�� 	l   
  via2  
ɸ k�   
  via2  Y� ��   
  via2  �\ :p   
  via2  C� 	l   
  via2  �4 @H   
  via2  �8 �0   
  via2  )�p !�(   
  via2  ;� !�(   
  via   �� ��   
  via2  �x j�   
  via3  #l\ &74   
  via2  �` T�   
  via2  *�� BD   
  via2  '}`  ��   
  via4  	�� T`   
  via2  �D �x   
  via3  4� #۰   
  via2  { �x   
  via4  E� &�x   
  via2  r� �   
  via2  7� |   
  via2  �4 ��   
  via2  �p ��   
  via2  � 	l   
  via2  	D D   
  via2  	�\ C�   
  via2  , %�(   
  via2  t !�(   
  via2  �$ ��   
  via2  wD ��   
  via2  'H ��   
  via2  �� -   
  via2  ~< �p   
  via2  �� �h   
  via2  	׈ Px   
  via2  5�    
  via2  $� �   
  via2  ��  �l   
  via2  r�  �l   
  via2  w�  ,�   
  via2  +�  �l   
  via2  �� ��   
  via2  � �   
  via2  $հ ��   
  via2  #d� ��   
  via2  (PP D   
  via2  M� �h   
  via2  	9T j�   
  via2  B� ��   
  via2  Y�  �l   
  via2  !�� ��   
  via2  �\ �   
  via2  �( �8   
  via2  � ��   
  via3  I� �   
  via2  U� 	l   
  via2  \4 k�   
  via2  5  9�   
  via2  %�� j�   
  via2  pp !�(   
  via2  4, gX   
  via2  &Ǽ P   
  via2  O� !�   
  via2  $H ��   
  via2  	�, &
H   
  via2  	�\ �   
  via2  "�| $I   
  via2  J� %�8   
  via2  "�L #��   
  via2   ?� #۰   
  via2  #��  �4   
  via2    �l   
  via2  ,�� @H   
  via2  H @H   
  via2  �� gX   
  via2  � @H   
  via2  )��    
  via2  '�� ��   
  via   �\ �   
  via2  ǜ #۰   
  via2  '�� �h   
  via2  Z� %�8   
  via2  D )h   
  via2  /D �0   
  via2  *� �x   
  via2  ,� ��   
  via3  � ��   
  via2  #ht �h   
  via2  #f� "�    
  via2  A� %�8   
  via   *�\    
  via2  "�� �   
  via2   .H ��   
  via2  (� ��   
  via2  �� @   
  via2  �$ �    
  via2  %8 ��   
  via2  -r� #۰   
  via2  -v� $�   
  via2  �l ]   
  via2  �8 9�   
  via2  �� 
�T   
  via2  #�8  �l   
  via2  !=� ��   
  via2  v�  �l   
  via3  )  @   
  via2  )�x �x   
  via2  %� �   
  via2  %�8 �   
  via2  0 %�8   
  via2  �� %�8   
  via2  &L� !�(   
  via2  (�x !�(   
  via2  �\ D   
  via2  2� T�   
  via2  :L �    
  via2  jL D   
  via2  ��     
  via2  ܌ D   
  via2  
b4 �x   
  via2  Ѩ �h   
  via2  #& #$   
  via2  o( j�   
  via2  )�l ��   
  via2  '�8 Al   
  via   )�  ʈ   
  via2  '�4 �x   
  via2  )�� �0   
  via3  %dD �x   
  via2  &d  �x   
  via2  "KL �h   
  via2  n� !�(   
  via2  �L �   
  via2  "j� 	!�   
  via2  '�4 	l   
  via2  "l �    
  via2  ,�� �0   
  via2   p� ��   
  via2  !�� j�   
  via2  �X $�`   
  via2  �� ��   
  via   p    
  via2  B` ��   
  via2   �  �4   
  via2  "=�  �l   
  via   > ��   
  via2  	7` @H   
  via2  �� �   
  via2  �� D   
  via3  E0 #��   
  via2  �4 !�(   
  via   m� $��   
  via2  !C� !�(   
  via2  +� �   
  via2  I` �   
  via2  N� ��   
  via2  f� ��   
  via2  *:� �   
  via2  &%� ��   
  via2  (� "`   
  via2  %�  #۰   
  via2  &� "d�   
  via2  $` #۰   
  via   `� ��   
  via2  C` j�   
  via2  T� C�   
  via2  �` D   
  via2  �X |�   
  via2  2� j�   
  via2  � �8   
  via2  )� �h   
  via2  (�� ~�   
  via2  %� !�(   
  via2  $� �   
  via2  W� �x   
  via2  $X� 9�   
  via2  �X �   
  via2  �t �   
  via2  �t 9�   
  via3  �� �   
  via2  �t ��   
  via2  ,ք �   
  via2  -�h ��   
  via2  �� %�8   
  via2  ~� %�8   
  via2  ,� o�   
  via2  %X�    
  via2  )d    
  via2  v� �h   
  via2  %5d C�   
  via2  �� x�   
  via2  ��  �l   
  via2  �P �h   
  via2  	�D �h   
  via2  �x k�   
  via2  �� 9�   
  via2  �l �   
  via2  �, �x   
  via2  !�d �   
  via2  �\  ��   
  via4  0� w�   
  via2  )@� ��   
  via2  )�� ��   
  via2  P �   
  via3  *a� �   
  via2  *:� #$   
  via2  �X Ը   
  via2  #�� �   
  via2  ,M� D   
  via2  -�, j�   
  via2  ,� �   
  via2  ,� #$   
  via2  + o�   
  via2  )P,     
  via2  -|� ��   
  via2  *� D   
  via2  '�    
  via2  "�h ��   
  via   wd �\   
  via2  *d �   
  via2  �  ��   
  via2  #�� �   
  via4  �L @   
  via2  -� ��   
  via3  )�H j�   
  via2  %X� j�   
  via2  #H ��   
  via2  )) D   
  via2  )�\ D   
  via2  +�� ��   
  via3  � %�8   
  via2  $-� �   
  via2  '�L g�   
  via2  28 #۰   
  via3  $�D �   
  via2  �� �x   
  via3  %Ѥ 9�   
  via2  �� 	l   
  via2  )d ��   
  via2  *X  �l   
  via2  &� Θ   
  via2  '�� D   
  via2  "߼ �l   
  via2  %}� Al   
  via3  -E� j�   
  via2  &� 9�   
  via2  �� h|   
  via2  c� Al   
  via2  Ȝ #۰   
  via2  !9� �   
  via2  �� �0   
  via2  ;� �X   
  via   	�� ��   
  via2  	9T Al   
  via2  $�D �    
  via2  '� ��   
  via2  )Dt $p    
  via2  -�t #۰   
  via2  +J ��   
  via2  %�� �0   
  via   2T '   
  via2  �D �h   
  via2  �p �   
  via2  �� 	l   
  via2  I� -   
  via2  V �h   
  via2   �0 	l   
  via2  X Al   
  via2  � -   
  via2  � �0   
  via2  %/� gX   
  via2  �\ @H   
  via2  "� ��   
  via2   %�8   
  via2  &�, �|   
  via2  V� Al   
  via2  $'� ��   
  via2  � �   
  via2  �4 %�(   
  via2  	�� !�(   
  via2  
=  ��   
  via2  <� %�8   
  via3    ,   
  via2  H� ��   
  via2  �� %�    
  via2  X #۰   
  via2  *ڴ @H   
  via2   $� 	l   
  via2  *� �    
  via2  )LD �0   
  via3  �� "��   
  via2  s� ��   
  via2  �L  �\   
  via2  �  �l   
  via2  /� �   
  via2  �D  �l   
  via2    D   
  via2  X Al   
  via4  	� ��   
  via2  4 9�   
  via2  4L �(   
  via2  R 9�   
  via2  *d �   
  via2  
�t D   
  via2  ^� D   
  via2  i� ��   
  via2  E, ��   
  via2  � ��   
  via2  `� `�   
  via2  ��  �l   
  via2  7�    
  via2  W�  �l   
  via2  �, ��   
  via2  	��  �l   
  via3  Ѩ  �<   
  via2  �D ��   
  via2  �� �   
  via2  �� 9�   
  via2  �� $��   
  via2  &� �   
  via2  ,\ �x   
  via2  f` @H   
  via2  �� %�8   
  via2  �4 !�(   
  via2  &74 `   
  via2  !�� 9�   
  via2    FL   
  via2  l ��   
  via2  ��  �\   
  via2  �� 9�   
  via   kd Sl   
  via2  A  	l   
  via2  �� 	l   
  via2  Ҡ �   
  via2  Ј ��   
  via2  ET %�8   
  via2  �H "h�   
  via2  ( �x   
  via2  �� #H   
  via2  t #۰   
  via   !tt  ʈ   
  via2  *�h !�(   
  via2  +�� f�   
  via2  "ph �0   
  via2  � �   
  via2  x� �   
  via2  &k�  �   
  via2  #jh #۰   
  via2  � �h   
  via2  f� �x   
  via3  +��    
  via2  ,�  �   
  via2  ,�� 9�   
  via2  � !�(   
  via2  ' ��   
  via2  � @H   
  via2  ;� !�8   
  via2  -�  �x   
  via2  .� �   
  via2  �( �0   
  via   !�� ]�   
  via2  !�  D   
  via2  "($ ��   
  via2  �� �   
  via3  � %�(   
  via2  (<� �   
  via2  4 �4   
  via2  �( Al   
  via2  � U�   
  via2  b� ��   
  via2  !, 8   
  via2  '!� ��   
  via2  �D k    
  via2  V� 	l   
  via2  Z� �h   
  via2  z4 �x   
  via2  #� 8   
  via2  5h �x   
  via2  -� Ј   
  via2     !�(   
  via2  +.� �   
  via2  -p �   
  via4  &�H �@   
  via2  �( @H   
  via3  $N� Θ   
  via2  	�( %�8   
  via2  %� "Ep   
  via2  �� !�(   
  via2  �� ��   
  via2  	H� ��   
  via4  .6 #۰   
  via2  ,�� #۰   
  via2  J %�    
  via2  m4 %�8   
  via   $V� 
�T   
  via2  g %�8   
  via2  	�� -   
  via2  � �h   
  via2  	�� �@   
  via2  �P �h   
  via   ut ��   
  via2  F� �   
  via2  � #CX   
  via2  "x %�8   
  via2  �d �   
  via2  �P �   
  via2  }      
  via2  �x j�   
  via   �� $   
  via2  � ��   
  via3  %ϰ �   
  via2  �( %�8   
  via3   �P %�(   
  via2  .t �0   
  via2  #�d 9�   
  via2  x ��   
  via2   �L �   
  via2  3� �   
  via2  +� %�@   
  via2  %�@ %�8   
  via2  (L  �\   
  via2  �8 	l   
  via2  � �   
  via2  j$ Al   
  via3  @H !�   
  via2  '7 �   
  via2  e$ ��   
  via2  K�  �l   
  via2  � $l8   
  via2  +�x D   
  via2  +� ��   
  via2  '� �   
  via2  �� Ј   
  via2  �� �   
  via2  -�H @H   
  via2  ,�� �x   
  via2  �� 4   
  via2  �� 9�   
  via2  (p ��   
  via2  #� 9�   
  via2  �� �h   
  via2   D ��   
  via2  � aX   
  via2  %�D !�(   
  via2  �4 �X   
  via2  }� �   
  via3  �P �   
  via2  �� �   
  via2  %�,  ܴ   
  via2  ؄ j�   
  via2  �� !��   
  via2  F !�(   
  via2  )�� ��   
  via2  (�� ��   
  via3  '�4 �\   
  via2  �� �x   
  via2  Q0 %�8   
  via2  .� D   
  via2  *il !�   
  via2  )�� !�(   
  via   	� 
�,   
  via2  � T�   
  via2  !�P %�8   
  via2  �� %�8   
  via3  �( 
�D   
  via2  &=  ��   
  via2  � 9�   
  via2  � ��   
  via2  "�8 x�   
  via2  � ��   
  via2  '� ��   
  via2  !�h ��   
  via2  �� j�   
  via2  �� #۰   
  via2  '� j�   
  via2  �� �h   
  via2  �( 
�   
  via2  �L ��   
  via2  
;$ �|   
  via2   Al   
  via2  
�X P   
  via2  V4 !�(   
  via2  �0 Al   
  via2  �� Al   
  via2  � !��   
  via2  �4 %�8   
  via2  �p !�(   
  via2  ,�� �h   
  via2  { ��   
  via2  "�l ��   
  via2  Wx �x   
  via2  ,�l j�   
  via2  �� �x   
  via2  $�l ��   
  via4  ��    
  via2  �� Al   
  via2  I� 
(   
  via2  �� �0   
  via2  d #��   
  via2  �� �   
  via  �  B�        �� ^� +  ,VR_NO_BUS    
  via    | l�   
  via    | ��   
  via2  3� �8   
  via2  .� �8   
  via2  �� �h   
  via2  	G  �h   
  via2  �L  ��   
  via3  .UT Ԙ   
  via   0� �   
  via   )� %)�   
  via2  )� %�8   
  via2  ,.� ��   
  via2  +v� D   
  via2  �0 %u�   
  via  �  B�        /� 6h +  ,VR_NO_BUS    
  via  �  B�        0� 6h +  ,VR_NO_BUS    
  via  �  B�        07� 6h +  ,VR_NO_BUS    
  via  �  B�        0^� 6h +  ,VR_NO_BUS    
  via  �  B�        /  .� +  ,VR_NO_BUS    
  via  �  B�         �� %)� +  ,VR_NO_BUS    
  via  �  B�         �� %)� +  ,VR_NO_BUS    
  via  �  B�        $� %)� +  ,VR_NO_BUS    
  via  �  B�        L %)� +  ,VR_NO_BUS    
  via  �  B�         �� #"$ +  ,VR_NO_BUS    
  via  �  B�        /� %)� +  ,VR_NO_BUS    
  via  �  B�        0� %)� +  ,VR_NO_BUS    
  via  �  B�        07� %)� +  ,VR_NO_BUS    
  via  �  B�        0^� %)� +  ,VR_NO_BUS    
  via  �  B�        / #"$ +  ,VR_NO_BUS    
  via  �  B�         ��  .� +  ,VR_NO_BUS    
  via  �  B�         ��  .� +  ,VR_NO_BUS    
  via  �  B�        $�  .� +  ,VR_NO_BUS    
  via  �  B�        L  .� +  ,VR_NO_BUS    
  via3  ('L ��   
  via  �  B�        /�  .� +  ,VR_NO_BUS    
  via  �  B�        0�  .� +  ,VR_NO_BUS    
  via  �  B�        07�  .� +  ,VR_NO_BUS    
  via  �  B�        0^�  .� +  ,VR_NO_BUS    
  via  �  B�         �� %)� +  ,VR_NO_BUS    
  via  �  B�         �� 6h +  ,VR_NO_BUS    
  via  �  B�         �� 6h +  ,VR_NO_BUS    
  via  �  B�        $� 6h +  ,VR_NO_BUS    
  via  �  B�        L 6h +  ,VR_NO_BUS    
  via  �  B�         ��  .� +  ,VR_NO_BUS    
  via  �  B�        /� B� +  ,VR_NO_BUS    
  via  �  B�        0� B� +  ,VR_NO_BUS    
  via  �  B�        07� B� +  ,VR_NO_BUS    
  via  �  B�        0^� B� +  ,VR_NO_BUS    
  via  �  B�        / 
�@ +  ,VR_NO_BUS    
  via  �  B�         �� !� +  ,VR_NO_BUS    
  via  �  B�         �� !� +  ,VR_NO_BUS    
  via  �  B�        $� !� +  ,VR_NO_BUS    
  via  �  B�        L !� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        /� !� +  ,VR_NO_BUS    
  via  �  B�        0� !� +  ,VR_NO_BUS    
  via  �  B�        07� !� +  ,VR_NO_BUS    
  via  �  B�        0^� !� +  ,VR_NO_BUS    
  via  �  B�        / �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        $� �� +  ,VR_NO_BUS    
  via  �  B�        L �� +  ,VR_NO_BUS    
  via  �  B�         �� �X +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        0� �� +  ,VR_NO_BUS    
  via  �  B�        07� �� +  ,VR_NO_BUS    
  via  �  B�        0^� �� +  ,VR_NO_BUS    
  via  �  B�        / �X +  ,VR_NO_BUS    
  via  �  B�         �� B� +  ,VR_NO_BUS    
  via  �  B�         �� B� +  ,VR_NO_BUS    
  via  �  B�        $� B� +  ,VR_NO_BUS    
  via  �  B�        L B� +  ,VR_NO_BUS    
  via  �  B�         �� 
�@ +  ,VR_NO_BUS    
  via  �  B�        /� � +  ,VR_NO_BUS    
  via  �  B�        0� � +  ,VR_NO_BUS    
  via  �  B�        07� � +  ,VR_NO_BUS    
  via  �  B�        0^� � +  ,VR_NO_BUS    
  via  �  B�        / �L +  ,VR_NO_BUS    
  via  �  B�         �� �X +  ,VR_NO_BUS    
  via  �  B�         �� �X +  ,VR_NO_BUS    
  via  �  B�        $� �X +  ,VR_NO_BUS    
  via  �  B�        L �X +  ,VR_NO_BUS    
  via  �  B�         �� 6h +  ,VR_NO_BUS    
  via  �  B�        /� �X +  ,VR_NO_BUS    
  via  �  B�        0� �X +  ,VR_NO_BUS    
  via  �  B�        07� �X +  ,VR_NO_BUS    
  via  �  B�        0^� �X +  ,VR_NO_BUS    
  via  �  B�        / 6h +  ,VR_NO_BUS    
  via  �  B�         �� 
�@ +  ,VR_NO_BUS    
  via  �  B�         �� 
�@ +  ,VR_NO_BUS    
  via  �  B�        $� 
�@ +  ,VR_NO_BUS    
  via  �  B�        L 
�@ +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        /� 
�@ +  ,VR_NO_BUS    
  via  �  B�        0� 
�@ +  ,VR_NO_BUS    
  via  �  B�        07� 
�@ +  ,VR_NO_BUS    
  via  �  B�        0^� 
�@ +  ,VR_NO_BUS    
  via  �  B�        / �� +  ,VR_NO_BUS    
  via  �  B�         �� � +  ,VR_NO_BUS    
  via  �  B�         �� � +  ,VR_NO_BUS    
  via  �  B�        $� � +  ,VR_NO_BUS    
  via  �  B�        L � +  ,VR_NO_BUS    
  via  �  B�         �� �L +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        0� �� +  ,VR_NO_BUS    
  via  �  B�        07� �� +  ,VR_NO_BUS    
  via  �  B�        0^� �� +  ,VR_NO_BUS    
  via  �  B�        / B� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        $� �� +  ,VR_NO_BUS    
  via  �  B�        L �� +  ,VR_NO_BUS    
  via  �  B�         �� � +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        0� �� +  ,VR_NO_BUS    
  via  �  B�        07� �� +  ,VR_NO_BUS    
  via  �  B�        0^� �� +  ,VR_NO_BUS    
  via  �  B�        / � +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        $� �� +  ,VR_NO_BUS    
  via  �  B�        L �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        0� �� +  ,VR_NO_BUS    
  via  �  B�        07� �� +  ,VR_NO_BUS    
  via  �  B�        0^� �� +  ,VR_NO_BUS    
  via  �  B�        / �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        $� �� +  ,VR_NO_BUS    
  via  �  B�        L �� +  ,VR_NO_BUS    
  via  �  B�         �� B� +  ,VR_NO_BUS    
  via  �  B�        /� �L +  ,VR_NO_BUS    
  via  �  B�        0� �L +  ,VR_NO_BUS    
  via  �  B�        07� �L +  ,VR_NO_BUS    
  via  �  B�        0^� �L +  ,VR_NO_BUS    
  via  �  B�        / �� +  ,VR_NO_BUS    
  via  �  B�         �� %� +  ,VR_NO_BUS    
  via  �  B�         �� %� +  ,VR_NO_BUS    
  via  �  B�        $� %� +  ,VR_NO_BUS    
  via  �  B�        L %� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        /� %� +  ,VR_NO_BUS    
  via  �  B�        0� %� +  ,VR_NO_BUS    
  via  �  B�        07� %� +  ,VR_NO_BUS    
  via  �  B�        0^� %� +  ,VR_NO_BUS    
  via  �  B�        / �� +  ,VR_NO_BUS    
  via  �  B�         �� Ll +  ,VR_NO_BUS    
  via  �  B�         �� Ll +  ,VR_NO_BUS    
  via  �  B�        $� Ll +  ,VR_NO_BUS    
  via  �  B�        L Ll +  ,VR_NO_BUS    
  via  �  B�         �� %� +  ,VR_NO_BUS    
  via  �  B�        /� Ll +  ,VR_NO_BUS    
  via  �  B�        0� Ll +  ,VR_NO_BUS    
  via  �  B�        07� Ll +  ,VR_NO_BUS    
  via  �  B�        0^� Ll +  ,VR_NO_BUS    
  via  �  B�        / %� +  ,VR_NO_BUS    
  via  �  B�         �� �L +  ,VR_NO_BUS    
  via  �  B�         �� �L +  ,VR_NO_BUS    
  via  �  B�        $� �L +  ,VR_NO_BUS    
  via  �  B�        L �L +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        /� #"$ +  ,VR_NO_BUS    
  via  �  B�        0� #"$ +  ,VR_NO_BUS    
  via  �  B�        07� #"$ +  ,VR_NO_BUS    
  via  �  B�        0^� #"$ +  ,VR_NO_BUS    
  via  �  B�        / !� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        $� �� +  ,VR_NO_BUS    
  via  �  B�        L �� +  ,VR_NO_BUS    
  via  �  B�         �� Ll +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        0� �� +  ,VR_NO_BUS    
  via  �  B�        07� �� +  ,VR_NO_BUS    
  via  �  B�        0^� �� +  ,VR_NO_BUS    
  via  �  B�        / Ll +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        $� �� +  ,VR_NO_BUS    
  via  �  B�        L �� +  ,VR_NO_BUS    
  via  �  B�         �� �� +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        0� �� +  ,VR_NO_BUS    
  via  �  B�        07� �� +  ,VR_NO_BUS    
  via  �  B�        0^� �� +  ,VR_NO_BUS    
  via  �  B�        / �� +  ,VR_NO_BUS    
  via  �  B�         �� #"$ +  ,VR_NO_BUS    
  via  �  B�         �� #"$ +  ,VR_NO_BUS    
  via  �  B�        $� #"$ +  ,VR_NO_BUS    
  via  �  B�        L #"$ +  ,VR_NO_BUS    
  via  �  B�         �� !� +  ,VR_NO_BUS    
  via  �  B�        /� &�\ +  ,VR_NO_BUS    
  via  �  B�        /=� &�\ +  ,VR_NO_BUS    
  via  �  B�        /d� &�\ +  ,VR_NO_BUS    
  via  �  B�        /�� &�\ +  ,VR_NO_BUS    
  via  �  B�        .� $�� +  ,VR_NO_BUS    
  via  �  B�        �� 84 +  ,VR_NO_BUS    
  via  �  B�        �� 84 +  ,VR_NO_BUS    
  via  �  B�        �� 84 +  ,VR_NO_BUS    
  via  �  B�        � 84 +  ,VR_NO_BUS    
  via  �  B�        �� �8 +  ,VR_NO_BUS    
  via  �  B�        /� 84 +  ,VR_NO_BUS    
  via  �  B�        /=� 84 +  ,VR_NO_BUS    
  via  �  B�        /d� 84 +  ,VR_NO_BUS    
  via  �  B�        /�� 84 +  ,VR_NO_BUS    
  via  �  B�        .� �8 +  ,VR_NO_BUS    
  via  �  B�        �� �T +  ,VR_NO_BUS    
  via  �  B�        �� �T +  ,VR_NO_BUS    
  via  �  B�        �� �T +  ,VR_NO_BUS    
  via  �  B�        � �T +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        /� �T +  ,VR_NO_BUS    
  via  �  B�        /=� �T +  ,VR_NO_BUS    
  via  �  B�        /d� �T +  ,VR_NO_BUS    
  via  �  B�        /�� �T +  ,VR_NO_BUS    
  via  �  B�        .� �� +  ,VR_NO_BUS    
  via  �  B�        �� &�\ +  ,VR_NO_BUS    
  via  �  B�        �� &�\ +  ,VR_NO_BUS    
  via  �  B�        �� &�\ +  ,VR_NO_BUS    
  via  �  B�        � &�\ +  ,VR_NO_BUS    
  via  �  B�        �� $�� +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        /=� �� +  ,VR_NO_BUS    
  via  �  B�        /d� �� +  ,VR_NO_BUS    
  via  �  B�        /�� �� +  ,VR_NO_BUS    
  via  �  B�        .� �� +  ,VR_NO_BUS    
  via  �  B�        �� 4l +  ,VR_NO_BUS    
  via  �  B�        �� 4l +  ,VR_NO_BUS    
  via  �  B�        �� 4l +  ,VR_NO_BUS    
  via  �  B�        � 4l +  ,VR_NO_BUS    
  via  �  B�        �� � +  ,VR_NO_BUS    
  via  �  B�        /� 4l +  ,VR_NO_BUS    
  via  �  B�        /=� 4l +  ,VR_NO_BUS    
  via  �  B�        /d� 4l +  ,VR_NO_BUS    
  via  �  B�        /�� 4l +  ,VR_NO_BUS    
  via  �  B�        .� � +  ,VR_NO_BUS    
  via  �  B�        �� � +  ,VR_NO_BUS    
  via  �  B�        �� � +  ,VR_NO_BUS    
  via  �  B�        �� � +  ,VR_NO_BUS    
  via  �  B�        � � +  ,VR_NO_BUS    
  via  �  B�        �� �T +  ,VR_NO_BUS    
  via  �  B�        /� � +  ,VR_NO_BUS    
  via  �  B�        /=� � +  ,VR_NO_BUS    
  via  �  B�        /d� � +  ,VR_NO_BUS    
  via  �  B�        /�� � +  ,VR_NO_BUS    
  via  �  B�        .� �T +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        � �� +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        /� �8 +  ,VR_NO_BUS    
  via  �  B�        /=� �8 +  ,VR_NO_BUS    
  via  �  B�        /d� �8 +  ,VR_NO_BUS    
  via  �  B�        /�� �8 +  ,VR_NO_BUS    
  via  �  B�        .� �� +  ,VR_NO_BUS    
  via  �  B�        �� 5� +  ,VR_NO_BUS    
  via  �  B�        �� 5� +  ,VR_NO_BUS    
  via  �  B�        �� 5� +  ,VR_NO_BUS    
  via  �  B�        � 5� +  ,VR_NO_BUS    
  via  �  B�        �� . +  ,VR_NO_BUS    
  via  �  B�        /� 5� +  ,VR_NO_BUS    
  via  �  B�        /=� 5� +  ,VR_NO_BUS    
  via  �  B�        /d� 5� +  ,VR_NO_BUS    
  via  �  B�        /�� 5� +  ,VR_NO_BUS    
  via  �  B�        .� . +  ,VR_NO_BUS    
  via  �  B�        �� ܐ +  ,VR_NO_BUS    
  via  �  B�        �� ܐ +  ,VR_NO_BUS    
  via  �  B�        �� ܐ +  ,VR_NO_BUS    
  via  �  B�        � ܐ +  ,VR_NO_BUS    
  via  �  B�        / %)� +  ,VR_NO_BUS    
  via  �  B�        /� ܐ +  ,VR_NO_BUS    
  via  �  B�        /=� ܐ +  ,VR_NO_BUS    
  via  �  B�        /d� ܐ +  ,VR_NO_BUS    
  via  �  B�        /�� ܐ +  ,VR_NO_BUS    
  via  �  B�        �� &�\ +  ,VR_NO_BUS    
  via  �  B�        �� �8 +  ,VR_NO_BUS    
  via  �  B�        �� �8 +  ,VR_NO_BUS    
  via  �  B�        �� �8 +  ,VR_NO_BUS    
  via  �  B�        � �8 +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        /�  �� +  ,VR_NO_BUS    
  via  �  B�        /=�  �� +  ,VR_NO_BUS    
  via  �  B�        /d�  �� +  ,VR_NO_BUS    
  via  �  B�        /��  �� +  ,VR_NO_BUS    
  via  �  B�        .� 4l +  ,VR_NO_BUS    
  via2  Z� "�    
  via  �  B�        �� ^� +  ,VR_NO_BUS    
  via  �  B�        �� ^� +  ,VR_NO_BUS    
  via  �  B�        � ^� +  ,VR_NO_BUS    
  via  �  B�        �� 84 +  ,VR_NO_BUS    
  via  �  B�        /� ^� +  ,VR_NO_BUS    
  via  �  B�        /=� ^� +  ,VR_NO_BUS    
  via  �  B�        /d� ^� +  ,VR_NO_BUS    
  via  �  B�        /�� ^� +  ,VR_NO_BUS    
  via  �  B�        .� 84 +  ,VR_NO_BUS    
  via  �  B�        �� "�L +  ,VR_NO_BUS    
  via  �  B�        �� "�L +  ,VR_NO_BUS    
  via  �  B�        �� "�L +  ,VR_NO_BUS    
  via  �  B�        � "�L +  ,VR_NO_BUS    
  via  �  B�        ��  �� +  ,VR_NO_BUS    
  via  �  B�        /� "�L +  ,VR_NO_BUS    
  via  �  B�        /=� "�L +  ,VR_NO_BUS    
  via  �  B�        /d� "�L +  ,VR_NO_BUS    
  via  �  B�        /�� "�L +  ,VR_NO_BUS    
  via  �  B�        .�  �� +  ,VR_NO_BUS    
  via  �  B�        ��  �� +  ,VR_NO_BUS    
  via  �  B�        ��  �� +  ,VR_NO_BUS    
  via  �  B�        ��  �� +  ,VR_NO_BUS    
  via  �  B�        �  �� +  ,VR_NO_BUS    
  via  �  B�        �� 4l +  ,VR_NO_BUS    
  via  �  B�        /� 
`@ +  ,VR_NO_BUS    
  via  �  B�        /=� 
`@ +  ,VR_NO_BUS    
  via  �  B�        /d� 
`@ +  ,VR_NO_BUS    
  via  �  B�        /�� 
`@ +  ,VR_NO_BUS    
  via  �  B�        .� 5� +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        � �� +  ,VR_NO_BUS    
  via  �  B�        �� ^� +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        /=� �� +  ,VR_NO_BUS    
  via  �  B�        /d� �� +  ,VR_NO_BUS    
  via  �  B�        /�� �� +  ,VR_NO_BUS    
  via  �  B�        .� ^� +  ,VR_NO_BUS    
  via  �  B�        �� . +  ,VR_NO_BUS    
  via  �  B�        �� . +  ,VR_NO_BUS    
  via  �  B�        �� . +  ,VR_NO_BUS    
  via  �  B�        � . +  ,VR_NO_BUS    
  via  �  B�        �� � +  ,VR_NO_BUS    
  via  �  B�        /� . +  ,VR_NO_BUS    
  via  �  B�        /=� . +  ,VR_NO_BUS    
  via  �  B�        /d� . +  ,VR_NO_BUS    
  via  �  B�        /�� . +  ,VR_NO_BUS    
  via  �  B�        .� � +  ,VR_NO_BUS    
  via  �  B�        �� 
`@ +  ,VR_NO_BUS    
  via  �  B�        �� 
`@ +  ,VR_NO_BUS    
  via  �  B�        �� 
`@ +  ,VR_NO_BUS    
  via  �  B�        � 
`@ +  ,VR_NO_BUS    
  via  �  B�        �� 5� +  ,VR_NO_BUS    
  via  �  B�        /� �� +  ,VR_NO_BUS    
  via  �  B�        /=� �� +  ,VR_NO_BUS    
  via  �  B�        /d� �� +  ,VR_NO_BUS    
  via  �  B�        /�� �� +  ,VR_NO_BUS    
  via  �  B�        .� 
`@ +  ,VR_NO_BUS    
  via  �  B�        �� $�� +  ,VR_NO_BUS    
  via  �  B�        �� $�� +  ,VR_NO_BUS    
  via  �  B�        �� $�� +  ,VR_NO_BUS    
  via  �  B�        � $�� +  ,VR_NO_BUS    
  via  �  B�        �� "�L +  ,VR_NO_BUS    
  via  �  B�        /� $�� +  ,VR_NO_BUS    
  via  �  B�        /=� $�� +  ,VR_NO_BUS    
  via  �  B�        /d� $�� +  ,VR_NO_BUS    
  via  �  B�        /�� $�� +  ,VR_NO_BUS    
  via  �  B�        .� "�L +  ,VR_NO_BUS    
  via  �  B�        �� � +  ,VR_NO_BUS    
  via  �  B�        �� � +  ,VR_NO_BUS    
  via  �  B�        �� � +  ,VR_NO_BUS    
  via  �  B�        � � +  ,VR_NO_BUS    
  via  �  B�        �� ܐ +  ,VR_NO_BUS    
  via  �  B�        /� � +  ,VR_NO_BUS    
  via  �  B�        /=� � +  ,VR_NO_BUS    
  via  �  B�        /d� � +  ,VR_NO_BUS    
  via  �  B�        /�� � +  ,VR_NO_BUS    
  via  �  B�        .� ܐ +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        �� �� +  ,VR_NO_BUS    
  via  �  B�        � �� +  ,VR_NO_BUS    
  via  �  B�        �� 
`@ +  ,VR_NO_BUS       !    , 0�@ 9� 1� 9� 1� Et 0�@ Et 0�@ 9�      !    , 0�@ ø 1� ø 1� �p 0�@ �p 0�@ ø      !    ,  � ��  @ ��  @ �D  � �D  � ��      !    , 0�@ �| 1� �| 1� �4 0�@ �4 0�@ �|      !    , 0�@ 't 1� 't 1� 3, 0�@ 3, 0�@ 't      !    ,  � %�\  @ %�\  @ %�  � %�  � %�\      !    , 0�@ �� 1� �� 1� �| 0�@ �| 0�@ ��      !    , 0�@ $ � 1� $ � 1� $� 0�@ $� 0�@ $ �      !    , 0�@  � 1�  � 1�   � 0�@   � 0�@  �      !    ,  � "�  @ "�  @ "߼  � "߼  � "�      !    , 0�@ 3t 1� 3t 1� ?, 0�@ ?, 0�@ 3t      !    , 0�@ �� 1� �� 1� �` 0�@ �` 0�@ ��      !    , 0�@ u� 1� u� 1� �L 0�@ �L 0�@ u�      !    , 0�@ i, 1� i, 1� t� 0�@ t� 0�@ i,      !    ,  � ��  @ ��  @ �`  � �`  � ��      !    , 0�@ � 1� � 1� �� 0�@ �� 0�@ �      !    ,  � {P  @ {P  @ �  � �  � {P      !    , 0�@  d 1�  d 1�  0�@  0�@  d      !    , 0�@ �< 1� �< 1� �� 0�@ �� 0�@ �<      !    ,  � &T  @ &T  @ &  � &  � &T      !    , 0�@ N� 1� N� 1� Z< 0�@ Z< 0�@ N�      !    , 0�@ �L 1� �L 1� � 0�@ � 0�@ �L      !    ,  � ֬  @ ֬  @ �d  � �d  � ֬      !    , 0�@ !0 1� !0 1� ,� 0�@ ,� 0�@ !0      !    ,  � N�  @ N�  @ Z<  � Z<  � N�      !    ,  � ��  @ ��  @ �T  � �T  � ��      !    ,  � !�\  @ !�\  @ "  � "  � !�\      !    ,  � d�  @ d�  @ p�  � p�  � d�      !    ,  � ��  @ ��  @ �d  � �d  � ��      !    ,  � ]�  @ ]�  @ iP  � iP  � ]�      !    , 0�@ �� 1� �� 1� �� 0�@ �� 0�@ ��      !    ,  � H  @ H  @ )   � )   � H      !    ,  � 7�  @ 7�  @ C�  � C�  � 7�      !    ,  � �   @ �   @ ��  � ��  � �       !    ,  � �  @ �  @ ��  � ��  � �      !    , 0�@ #�� 1� #�� 1� #� 0�@ #� 0�@ #��      !    ,  � ��  @ ��  @ ��  � ��  � ��      !    , 0�@ �| 1� �| 1� �4 0�@ �4 0�@ �|      !    , 0�@ � 1� � 1� d 0�@ d 0�@ �      !    , 0�@ � 1� � 1� � 0�@ � 0�@ �      !    , 0�@ �� 1� �� 1� � 0�@ � 0�@ ��          , �x &� �0 &� �0 '< �x '< �x &�          , ,��     -@     -@  � ,��  � ,��              , -i      -t�     -t�  � -i   � -i               , *��     *�8     *�8  � *��  � *��              , .$�     .08     .08  � .$�  � .$�              , *<�     *H8     *H8  � *<�  � *<�              ,  x�      �8      �8  �  x�  �  x�              ,  20      =�      =�  �  20  �  20              , &5@     &@�     &@�  � &5@  � &5@              , )��     )�     )�  � )��  � )��              , )�X     )�     )�  � )�X  � )�X              , (!p     (-(     (-(  � (!p  � (!p              , � &� �� &� �� '< � '< � &�          , � &� �� &� �� '< � '< � &�          , 8� &� D� &� D� '< 8� '< 8� &�          , %��     %ϰ     %ϰ  � %��  � %��              , �L &� � &� � '< �L '< �L &�          , ;� &� G� &� G� '< ;� '< ;� &�          , �H     �      �   � �H  � �H              , $�p &� $�( &� $�( '< $�p '< $�p &�          , &��     &ό     &ό  � &��  � &��              , $X�     $dh     $dh  � $X�  � $X�              , u( &� �� &� �� '< u( '< u( &�          , e� &� q� &� q� '< e� '< e� &�          , � &� �� &� �� '< � '< � &�          , H� &� T` &� T` '< H� '< H� &�          , .Ox     .[0     .[0  � .Ox  � .Ox              , $�(     $��     $��  � $�(  � $�(              , � &� �� &� �� '< � '< � &�          , 
͠     
�X     
�X  � 
͠  � 
͠              , %%� &� %1| &� %1| '< %%� '< %%� &�          , �p     (     (  � �p  � �p              , V�     b�     b�  � V�  � V�              , Rp     ^(     ^(  � Rp  � Rp              ,  d� &�  p� &�  p� '<  d� '<  d� &�          , #?p &� #K( &� #K( '< #?p '< #?p &�          , #r8 &� #}� &� #}� '< #r8 '< #r8 &�          , �� &� �p &� �p '< �� '< �� &�          , &4 &� 1� &� 1� '< &4 '< &4 &�          , 	�� &� 	�� &� 	�� '< 	�� '< 	�� &�          , 	E &� 	P� &� 	P� '< 	E '< 	E &�          , I &� T� &� T� '< I '< I &�          , � &� p &� p '< � '< � &�      1    ,  � �  @ �  @ I\  � I\  � �      1    , 0�@ �L 1� �L 1� n� 0�@ n� 0�@ �L      !    , $5� �L ,�d �L ,�d � $5� � $5� �L      !    , ,� 't 0� 't 0� 3, ,� 3, ,� 't      !    , � � 0� � 0� d � d � �      !    , �p  d 0�  d 0�  �p  �p  d      !    , )D �� "�� �� "�� �t )D �t )D ��      !    ,  d "� � "� � "߼  d "߼  d "�      !    , � &�� �� &�� �� 'T � 'T � &��      !    ,  d ֬  D\ ֬  D\ �d  d �d  d ֬      !    , � N< Z� N< Z� Y� � Y� � N<      !    , 	!�  N  ��  N  ��  Y� 	!�  Y� 	!�  N       !    , �  N  ��  N  ��  Y� �  Y� �  N       !    , ,*� N� 0� N� 0� Z< ,*� Z< ,*� N�      !    , $� @ )B� @ )B� � $� � $� @      !    ,  d 7� � 7� � C�  d C�  d 7�      !    ,  d &T  :� &T  :� &  d &  d &T      !    , %;@ _d &�� _d &�� k %;@ k %;@ _d      !    , &ɰ � '�H � '�H � &ɰ � &ɰ �      !    ,  d �� ?� �� ?� ��  d ��  d ��      !    ,  d �� |� �� |� �D  d �D  d ��      !    ,  � !�\ � !�\ � "  � "  � !�\      !    , �� !�� T` !�� T` !�d �� !�d �� !��      !    , ,�� �� 0� �� 0� �� ,�� �� ,�� ��      !    , �� #T �� #T �� #& �� #& �� #T      !    ,  d {P _H {P _H �  d �  d {P      !    , �� &l X� &l X� &$ �� &$ �� &l      !    ,  d %�\ � %�\ � %�  d %�  d %�\      !    ,  �� s� �� s� �l  �l  ��      !    , &�l �d 0�� �d 0�� � &�l � &�l �d      !    , u� j$ �  j$ �  u� u� u� u� j$      !    ,  � S� *� S� *� _�  � _�  � S�      !    , ؀ !�� �@ !�� �@ !� ؀ !� ؀ !��      !    , 4, q� �4 q� �4 }d 4, }d 4, q�      !    , ,�p �L 0� �L 0� � ,�p � ,�p �L      !    , /h &+| " T &+| " T &74 /h &74 /h &+|      !    , 	H� &�� 	w� &�� 	w� 'T 	H� 'T 	H� &��      !    , #Ad #�� $�  #�� $�  $� #Ad $� #Ad #��      !    , ,�� � -n� � -n� �� ,�� �� ,�� �      !    , p� a| &R� a| &R� m4 p� m4 p� a|      !    , v� �� �� �� �� �t v� �t v� ��      !    ,  d � 
� � 
� ��  d ��  d �      !    , W� �� !�d �� !�d ۴ W� ۴ W� ��      !    , �4 &�� � &�� � 'T �4 'T �4 &��      !    , � H� � H� � T@ � T@ � H�      !    , )� �� *(� �� *(� �P )� �P )� ��      !    , �` �L !�� �L !�� � �` � �` �L      !    ,  �� 
�� $�� 
�� $�� P  �� P  �� 
��      !    ,  d N� �  N� �  Z<  d Z<  d N�      !    , 
� 	� d  	� d  X 
� X 
� 	�      !    , (, eh �� eh �� q  (, q  (, eh      !    , 	�� &�� 	Ք &�� 	Ք 'T 	�� 'T 	�� &��      !    , ?� &�� n� &�� n� 'T ?� 'T ?� &��      !    , �( �� *:� �� *:� �x �( �x �( ��      !    , � � _� � _� �p � �p � �      !    , $l8 1� '�� 1� '�� =� $l8 =� $l8 1�      !    , $�H :� *d :� *d Fp $�H Fp $�H :�      !    , %Ә 9� 0� 9� 0� Et %Ә Et %Ә 9�      !    , #H "l *�l "l *�l "($ #H "($ #H "l      !    , 
 !9� �l !9� �l !E� 
 !E� 
 !9�      !    , �� �� �� �� �� �� �� �� �� ��      !    , �4 	D p� 	D p� 	� �4 	� �4 	D      !    , 
Zd DX � DX � P 
Zd P 
Zd DX      !    , '� qd V� qd V� } '� } '� qd      !    , )y0 d� ."� d� ."� pL )y0 pL )y0 d�      !    , -c$ �< 0� �< 0� �� -c$ �� -c$ �<      !    , *�( �� 0� �� 0� �` *�( �` *�( ��      !    , n0 :l cp :l cp F$ n0 F$ n0 :l      !    , I� � �x � �x �L I� �L I� �      !    , &� & � �� & � �� &< &� &< &� & �      !    , 
;$ 	�` {P 	�` {P 	� 
;$ 	� 
;$ 	�`      !    , �H 
͠ �` 
͠ �` 
�X �H 
�X �H 
͠      !    , �� &�� �� &�� �� 'T �� 'T �� &��      !    , !�� �� &�� �� &�� �� !�� �� !�� ��      !    , � N� 
 � N� 
 � Z< � Z< � N�      !    , �x C\ S� C\ S� O �x O �x C\      !    , �� �� �� �� �� �� �� �� �� ��      !    , #z  ' '�d  ' '�d  2� #z  2� #z  '      !    , �� �  M  �  M  �� �� �� �� �       !    ,  d �� �� �� �� �d  d �d  d ��      !    , �� 
͠ _  
͠ _  
�X �� 
�X �� 
͠      !    , � D $� D $� "� � "� � D      !    , , "�, 	;H "�, 	;H #� , #� , "�,      !    , :p �� iP �� iP �� :p �� :p ��      !    , ~� 
�� � 
�� � 
�� ~� 
�� ~� 
��      !    , "�(  � 0�  � 0�   � "�(   � "�(  �      !    , 'o� � 0� � 0� �� 'o� �� 'o� �      !    , �T 3� F( 3� F( ?x �T ?x �T 3�      !    , �� 	;H 
j 	;H 
j 	G  �� 	G  �� 	;H      !    , ݈ H �, H �, )  ݈ )  ݈ H      !    , *Q� !0 0� !0 0� ,� *Q� ,� *Q� !0      !    , $0 DX *]� DX *]� P $0 P $0 DX      !    , �� �� * �� * Ǡ �� Ǡ �� ��      !    , 'g� �� 0� �� 0� � 'g� � 'g� ��      !    , �� $פ )  $פ )  $�\ �� $�\ �� $פ      !    , ""H � -A� � -A� �t ""H �t ""H �      !    , *@ \� *gx \� *gx hX *@ hX *@ \�      !    ,  d �  �� �  �� ��  d ��  d �       !    , #?p &Xh #r8 &Xh #r8 &d  #?p &d  #?p &Xh      !    ,   �  � *�  *�        !    , q� &N� �� &N� �� &Z\ q� &Z\ q� &N�      !    , 'w�  � )�  � )�  �� 'w�  �� 'w�  �      !    , $�p '� $�8 '� $�8 '%| $�p '%| $�p '�      !    , �� 	� #�� 	� #�� X �� X �� 	�      !    , &T �P *k` �P *k` � &T � &T �P      !    , $հ &�� %-� &�� %-� 'T $հ 'T $հ &��      !    , 3, � �d � �d �� 3, �� 3, �      !    , #nP &�� #�0 &�� #�0 'T #nP 'T #nP &��      !    , #� �� �8 �� �8 Δ #� Δ #� ��      !    ,  d d� �D d� �D p�  d p�  d d�      !    , `� %=4 �� %=4 �� %H� `� %H� `� %=4      !    , DT �� � �� � �� DT �� DT ��      !    ,  d ]� � ]� � iP  d iP  d ]�      !    , )} �p +�8 �p +�8 �( )} �( )} �p      !    , .S` #�� 0�� #�� 0�� $� .S` $� .S` #��      !    , % �� �� �� �� �� % �� % ��      !    , T� % �� % �� %%� T� %%� T� %      !    , -T YH � YH � e  -T e  -T YH      !    , t� @ �� @ �� � t� � t� @      !    , 
� �  � �  � �p 
� �p 
� �      !    , .08 #�� 0� #�� 0� #� .08 #� .08 #��      !    , &  �� &�   �� &�   �x &  �x &  ��      !    , 	j( �\ W� �\ W� � 	j( � 	j( �\      !    , -�� #�� .;� #�� .;� $� -�� $� -�� #��      !    , 0� 	 �� 	 �� 	'� 0� 	'� 0� 	      !    , (�� 9x ,�( 9x ,�( E0 (�� E0 (�� 9x      !    , ,.� ø 0� ø 0� �p ,.� �p ,.� ø      !    , [  N  ׄ  N  ׄ  Y� [  Y� [  N       !    ,  .� &+| ~ &+| ~ &74  .� &74  .� &+|          , �  N  ��  N  �� X � X �  N           , ~� 
͠ �` 
͠ �` 
�� ~� 
�� ~� 
͠          , .$� �  .08 �  .08 �| .$� �| .$� �           , , "� '� "� '� #� , #� , "�          , � $�� �� $�� �� 'T � 'T � $��          , �D @l �� @l �� a4 �D a4 �D @l          , y4 6< �� 6< �� 'T y4 'T y4 6<          , 0�( �� 1� �� 1� "� 0�( "� 0�( ��          ,  � B�  � B�  � _�  � _�  � B�          , ,�� �� ,�x �� ,�x �T ,�� �T ,�� ��          , 9P 0� E 0� E "nt 9P "nt 9P 0�          , b� c� n� c� n� 'T b� 'T b� c�          , �X 	  	  �� �X �� �X 	          , �8 %$ �� %$ �� %H� �8 %H� �8 %$          , � & � �� & � �� &3L � &3L � & �          , "� &l " T &l " T &74 "� &74 "� &l          , ,��  � -@  � -@ �� ,�� �� ,��  �          , -e �� -p� �� -p� � -e � -e ��          , "�x !x "�0 !x "�0 !�� "�x !�� "�x !x          , �  ' ��  ' ��  Y� �  Y� �  '          , *@ �  *(� �  *(� � *@ � *@ �           , **� = *6� = *6� �� **� �� **� =          , %` �L % �L % �t %` �t %` �L          , 8� #�� D� #�� D� &� 8� &� 8� #��          , �x L �0 L �0 O �x O �x L          , "�x #�� "�0 #�� "�0 $N� "�x $N� "�x #��          , � ?t �� ?t �� �T � �T � ?t          , � N< X N< X  � �  � � N<          , N� z� Z� z� Z� Y� N� Y� N� z�          , &�x = '0 = '0 Rl &�x Rl &�x =          , �( % �� % �� &3L �( &3L �( %          , $�h #�� $�  #�� $�  $� $�h $� $�h #��          , #Ad #�� #M #�� #M $� #Ad $� #Ad #��          , rd &l ~ &l ~ &74 rd &74 rd &l          ,  .� &T  :� &T  :� &74  .� &74  .� &T          , ${� 
ш $�� 
ш $�� P ${� P ${� 
ш          , �H � �  � �  l �H l �H �          , �P $Ӽ � $Ӽ � &$ �P &$ �P $Ӽ          , $�T :l $� :l $� �\ $�T �\ $�T :l          , h "� #  "� #  $�d h $�d h "�          , #�h μ #�  μ #�  F$ #�h F$ #�h μ          , .Ox  � .[0  � .[0 �t .Ox �t .Ox  �          , *.� v� *:� v� *:� t� *.� t� *.� v�          , �� �� �h �� �h �� �� �� �� ��          , �( e� �� e� �� �x �( �x �( e�          , #b� � #nP � #nP �d #b� �d #b� �          , �� =� �h =� �h � �� � �� =�          , �� � �x � �x ?� �� ?� �� �          , 	l !$` 	w� !$` 	w� 'T 	l 'T 	l !$`          , �P �8 � �8 � p� �P p� �P �8          , 4, q� ?� q� ?� �� 4, �� 4, q�          , �H  � �   � �  �4 �H �4 �H  �          , 'o� � '{l � '{l �� 'o� �� 'o� �          , .S` #�� ._ #�� ._ $+� .S` $+� .S` #��          , � �� �� �� ��  Ơ �  Ơ � ��          , �L H � H � P �L P �L H          , 
Zd �8 
f �8 
f P 
Zd P 
Zd �8          , &'� ~@ &3L ~@ &3L 
)� &'� 
)� &'� ~@          , y4 �T �� �T �� /D y4 /D y4 �T          , 0�( �� 1� �� 1� �� 0�( �� 0�( ��          , H� !�L T` !�L T` &� H� &� H� !�L          ,  �D Đ  �� Đ  �� nX  �D nX  �D Đ          , �\ �� � �� � 'T �\ 'T �\ ��          , � �� �� �� �� !� � !� � ��          ,  �� 
ш  �x 
ш  �x P  �� P  �� 
ш          , & �x &� �x &� ?� & ?� & �x          , "�4 r� "�� r� "�� �t "�4 �t "�4 r�          , /  !Kp :� !Kp :� #� /  #� /  !Kp          , *�� � *�H � *�H �@ *�� �@ *�� �          , '� �� '�H �� '�H � '� � '� ��          , ({H � (�  � (�  2� ({H 2� ({H �          , R( �� ]� �� ]� �T R( �T R( ��          , �< "� �� "� �� $�t �< $�t �< "�          , ƀ ~� �8 ~� �8 Δ ƀ Δ ƀ ~�          , !�� �� !�� �� !�� ?� !�� ?� !�� ��          , #7� �� #CX �� #CX �H #7� �H #7� ��          , *� >4 *d >4 *d �t *� �t *� >4          , X� �D dH �D dH ( X� ( X� �D          , i d� t� d� t� �� i �� i d�          , *_� �P *k` �P *k` � *_� � *_� �P          , ,k n� ,v� n� ,v� �< ,k �< ,k n�          , E� Z� QP Z� QP 
� E� 
� E� Z�          , Sh 
͠ _  
͠ _  �� Sh �� Sh 
͠          , '� �$ '�� �$ '�� � '� � '� �$          , ~� �� �� �� �� �t ~� �t ~� ��          , *�@ �� *�� �� *�� /D *�@ /D *�@ ��          , �4 	D �� 	D �� 	� �4 	� �4 	D          , WT a| c a| c ڔ WT ڔ WT a|          , V�  � b�  � b�  �8 V�  �8 V�  �          , �� $�| 	� $�| 	� $�\ �� $�\ �� $�|          , &ɰ � &�h � &�h �� &ɰ �� &ɰ �          ,  �t 	� !, 	� !, F$  �t F$  �t 	�          , � �� � �� �  � �  � � ��          , 3, � >� � >� � 3, � 3, �          , (�p = (�( = (�( �� (�p �� (�p =          , \ 4 g� 4 g�   \   \ 4          , 
� �� 
'� �� 
'� %� 
� %� 
� ��          , ��  ' ��  ' ��  Y� ��  Y� ��  '          , \� :l h� :l h� "KL \� "KL \� :l          , �� "� �p "� �p &� �� &� �� "�          , �` `< � `< � � �` � �` `<          , I� � U� � U� � I� � I� �          , 	�� N� 
 � N� 
 � �L 	�� �L 	�� N�          , &ό eD &�D eD &�D � &ό � &ό eD          , �0 [ �� [ �� "�� �0 "�� �0 [          , %�p �8 %�( �8 %�( <d %�p <d %�p �8          , *��  � *�8  � *�8 ?� *�� ?� *��  �          , ,*� � ,6\ � ,6\ Px ,*� Px ,*� �          ,  � c�  X c�  X �x  � �x  � c�          , )} �p )�� �p )�� ,8 )} ,8 )} �p          , 'Pt �� '\, �� '\, k� 'Pt k� 'Pt ��          , ;  O� F� O� F� �� ;  �� ;  O�          , �� :l �� :l �� m4 �� m4 �� :l          , %;@ _d %F� _d %F� �d %;@ �d %;@ _d          , P 't ( 't ( �d P �d P 't          , XH  � d   � d  X XH X XH  �          , �� i� �@ i� �@ Ǡ �� Ǡ �� i�          , d �� * �� * Ǡ d Ǡ d ��          , - � �P -,t �P -,t f� - � f� - � �P          , � �� �� �� �� �L � �L � ��          , %�� 	׈ & � 	׈ & � y4 %�� y4 %�� 	׈          , ~� �� �� �� �� "($ ~� "($ ~� ��          , !�l b� !�$ b� !�$ � !�l � !�l b�          , �� !�� �@ !�� �@ !� �� !� �� !��          , +� :l 7� :l 7� �\ +� �\ +� :l          , )D r� 4� r� 4� �t )D �t )D r�          ,  20  �  =�  �  =� 	�0  20 	�0  20  �          , � !9� �l !9� �l !l� � !l� � !9�          , �( %�$ �� %�$ �� %� �( %� �( %�$          , &T �P & �P & GH &T GH &T �P          , -� d� -�� d� -�� � -� � -� d�          , �p � �( � �( g4 �p g4 �p �          , *@ �� 5� �� 5� �� *@ �� *@ ��          , �h !� �  !� �  #� �h #� �h !�          , �P #�� � #�� � $u� �P $u� �P #��          , 0� �� <� �� <� 	'� 0� 	'� 0� ��          , }h G� �  G� �  �� }h �� }h G�          , �� �( �� �( �� � �� � �� �(          , *@ �\ *(� �\ *(� ^� *@ ^� *@ �\          , ,� �D ,�� �D ,�� 3, ,� 3, ,� �D          , -� ET -�d ET -�d 	u� -� 	u� -� ET          , �� 	 �� 	 �� 	q� �� 	q� �� 	          , �� l< �p l< �p �D �� �D �� l<          , F� d� RL d� RL �| F� �| F� d�          , t� @ �x @ �x @ t� @ t� @          , $�D m| $�� m| $�� �� $�D �� $�D m|          , >x 0� J0 0� J0 �� >x �� >x 0�          , -i   � -t�  � -t� � -i  � -i   �          ,  i� � i� � L(  L(  i�          , #� �� /� �� /� �� #� �� #� ��          , �� = �� = �� &�l �� &�l �� =          , z| q� �4 q� �4 F$ z| F$ z| q�          , �, �, �� �, �� �� �, �� �, �,          , ̀ !�\ �8 !�\ �8 $� ̀ $� ̀ !�\          , � ٜ "P ٜ "P � � � � ٜ          , +� 7� +�� 7� +��  +�  +� 7�          , 	�  �8 	�� �8 	�� �� 	�  �� 	�  �8          , AD $�� L� $�� L� &�l AD &�l AD $��          , � !� �� !� �� "$< � "$< � !�          , ,*� N� ,6\ N� ,6\ �| ,*� �| ,*� N�          , &F� �P &R� �P &R� '0 &F� '0 &F� �P          , �< 
ɸ � 
ɸ � 
�� �< 
�� �< 
ɸ          , �H 
͠ �  
͠ �  �� �H �� �H 
͠          , @ �T � �T �  � @  � @ �T          , )� _� *� _� *� �P )� �P )� _�          , �� � �x � �x %\ �� %\ �� �          , �   @   @ 2� � 2� �            , �p  � (  � ( X �p X �p  �          , 
� 4 
�� 4 
�� �p 
� �p 
� 4          ,  d ��  % ��  % �T  d �T  d ��          ,  8� :l  D\ :l  D\ �d  8� �d  8� :l          , K qd V� qd V� $�< K $�< K qd          , � �� p �� p &� � &� � ��          , �� [ � [ � �� �� �� �� [          , � � 'T � 'T � � � � �          , !  �X ,�  �X ,�  �` !  �` !  �X          , �p  � �(  � �( b� �p b� �p  �          , 
;$ 	f@ 
F� 	f@ 
F� 	� 
;$ 	� 
;$ 	f@          , 
 %�$ 
!� %�$ 
!� %� 
 %� 
 %�$          , (� �4 (�� �4 (�� � (� � (� �4          , $0 H $%� H $%� P $0 P $0 H          , *Q� !0 *]� !0 *]� P *Q� P *Q� !0          , � �d (� �d (� /D � /D � �d          , ʌ d� �D d� �D �� ʌ �� ʌ d�          , ��  �  � _� �� _� ��           , Ј �T �@ �T �@ �t Ј �t Ј �T          , 	4 "�� � "�� � "߼ 	4 "߼ 	4 "��          , $� �� 0h �� 0h #ݤ $� #ݤ $� ��          ,  [4 :l  f� :l  f� &�l  [4 &�l  [4 :l          , � !8 �d !8 �d %� � %� � !8          , &4 "�� 1� "�� 1� &� &4 &� &4 "��          , U8 �� `� �� `� )  U8 )  U8 ��          , (, >X 3� >X 3� q  (, q  (, >X          , �� �� 	x �� 	x �� �� �� �� ��          , )��  � )�  � )�  @t )��  @t )��  �          , *�( �� *�� �� *�� 2� *�( 2� *�( ��          , #H �� #(  �� #(   � #H  � #H ��          , ""H x� ".  x� ".  �t ""H �t ""H x�          , -68 ʬ -A� ʬ -A� �t -68 �t -68 ʬ          , "�� D� "� D� "� �� "�� �� "�� D�          , %�` �h %� �h %� �� %�` �� %�` �h          , M� �| Y� �| Y�  M�  M� �|          , &�p 	�� &�( 	�� &�( �D &�p �D &�p 	��          , -?� � -K� � -K� p� -?� p� -?� �          , DT �� P �� P 	� DT 	� DT ��          , Qt x ], x ], /D Qt /D Qt x          , Xl H d$ H d$ G� Xl G� Xl H          , � �P X �P X 2� � 2� � �P          , &��  � ' `  � ' `  8 &��  8 &��  �          , ,�@ �� ,�� �� ,�� �� ,�@ �� ,�@ ��          , *ܨ �� *�` �� *�` �| *ܨ �| *ܨ ��          , 	�H 6� 	�  6� 	�  �T 	�H �T 	�H 6�          , s� Ҥ 8 Ҥ 8 � s� � s� Ҥ          , % � %#� � %#� �� % �� % �          , $�(  � $��  � $�� eH $�( eH $�(  �          , 
 !�4 � !�4 � " 
 " 
 !�4          , !�@ `< !�� `< !�� � !�@ � !�@ `<          , #?p &Xh #K( &Xh #K( &� #?p &� #?p &Xh          , W� :l cp :l cp m4 W� m4 W� :l          , +� ?t +p ?t +p 2� +� 2� +� ?t          , -�� #� -�h #� -�h �� -�� �� -�� #�          , #z  ' #��  ' #��  �H #z  �H #z  '          , +� � +d � +d �� +� �� +� �          , � �| *� �| *� �t � �t � �|          , #nP �� #z �� #z m #nP m #nP ��          , �t �( �, �( �, )  �t )  �t �(          , C� 	�� O` 	�� O` �� C� �� C� 	��          , �� �� 	� �� 	� 8| �� 8| �� ��          , %^h `< %j  `< %j  �T %^h �T %^h `<          , @  !�\ K� !�\ K� & @  & @  !�\          ,  �� 	�x  �| 	�x  �| K,  �� K,  �� 	�x          , �d 't  't  F$ �d F$ �d 't          , #�x ʬ #�0 ʬ #�0 'T #�x 'T #�x ʬ          , )�l 	�� )�$ 	�� )�$ pl )�l pl )�l 	��          , Z� 4 fd 4 fd �� Z� �� Z� 4          , �� �� �H �� �H �� �� �� �� ��          , "�� d� "�p d� "�p �t "�� �t "�� d�          , �� d� �� d� �� j� �� j� �� d�          , D � � � � iL D iL D �          , �  �� � �� � �D �  �D �  ��          , Ah �  M  �  M  )  Ah )  Ah �           ,  �� �h  �< �h  �< 
�@  �� 
�@  �� �h          , � � �� � �� �� � �� � �          , v� $�� �p $�� �p %�� v� %�� v� $��          , *.� �� *:� �� *:� x� *.� x� *.� ��          , !�p x !�( x !�( _� !�p _� !�p x          , �� �� �� �� �� )  �� )  �� ��          , +� �  7� �  7� �t +� �t +� �           , H m|   m|   #� H #� H m|          , ?t �� K, �� K, 	� ?t 	� ?t ��          , �� !=� �� !=� �� "nt �� "nt �� !=�          , u� C �p C �p u� u� u� u� C          , �� !�, 	� !�, 	� $�L �� $�L �� !�,          , 
 |� � |� � !� 
 !� 
 |�          , �D ?x �� ?x �� fd �D fd �D ?x          ,  �L D0  � D0  � �L  �L �L  �L D0          , %��  � %ϰ  � %ϰ c0 %�� c0 %��  �          , $� �0 $�� �0 $�� � $� � $� �0          , )6� �0 )B� �0 )B� � )6� � )6� �0          , �X 	f@  	f@  	� �X 	� �X 	f@          , v� ', �� ', �� m4 v� m4 v� ',          , p� :l |� :l |� m4 p� m4 p� :l          , 0�( �� 1� �� 1� ڔ 0�( ڔ 0�( ��          , �� !� ހ !� ހ !�d �� !�d �� !�          , ݈ �8 �@ �8 �@ )  ݈ )  ݈ �8          ,  x�  �  �8  �  �8 �   x� �   x�  �          , 7� 4 C� 4 C� jL 7� jL 7� 4          , -T 28 9 28 9 e  -T e  -T 28          ,  ��  � ��  � p�  p�  ��          , �� %�\ �P %�\ �P &$ �� &$ �� %�\          , 
�� �4 
�l �4 
�l 
H� 
�� 
H� 
�� �4          , �� � �P � �P p� �� p� �� �          , '� C 3� C 3� } '� } '� C          ,  �  � �  � 	q�  	q�  �          , � !�\ �� !�\ �� 'T � 'T � !�\          , �� #�� � #�� � %�� �� %�� �� #��          , �� 	�P ܌ 	�P ܌ 
H� �� 
H� �� 	�P          , H@ 
= S� 
= S� ø H@ ø H@ 
=          , &� & � 2X & � 2X &3L &� &3L &� & �          , `� %$ l< %$ l< %H� `� %H� `� %$          , �� 	j( ݨ 	j( ݨ 	�@ �� 	�@ �� 	j(          , &� �� &�� �� &�� А &� А &� ��          , �H j$ �  j$ �  /D �H /D �H j$          , DT ;� P ;� P �� DT �� DT ;�          , -|� P -�@ P -�@ s� -|� s� -|� P          , :p �� F( �� F( �� :p �� :p ��          , %�� � %Ռ � %Ռ Et %�� Et %�� �          , M  %�\ X� %�\ X� &$ M  &$ M  %�\          , 
}� 
�� 
�D 
�� 
�D � 
}� � 
}� 
��          , q  �� |� �� |� �T q  �T q  ��          , �P �< � �< � y| �P y| �P �<          , h �� s� �� s� �| h �| h ��          ,  �� *� �� *� �d  �d  ��          , Ќ !� �D !� �D " Ќ " Ќ !�          , W� � cP � cP �� W� �� W� �          , Lp �� X( �� X( �� Lp �� Lp ��          , �� �� �D �� �D �D �� �D �� ��          , � �l 	� �l 	� H� � H� � �l          , � �� 	� �� 	� �` � �` � ��          , �� !$` � !$` � #� �� #� �� !$`          , M�  �X Y�  �X Y� X M� X M�  �X          , �P g� � g� � �, �P �, �P g�          , ��  N  ׄ  N  ׄ  � ��  � ��  N           , [  ' f�  ' f�  Y� [  Y� [  '          , y � �� � �� C� y C� y �          , �P 28 � 28 � e  �P e  �P 28          , #�0  � #��  � #�� X #�0 X #�0  �          ,  8 ^�  � ^�  � 
  8 
  8 ^�          , s4 	f@ ~� 	f@ ~� 	� s4 	� s4 	f@          , �� 
͠ �� 
͠ �� ø �� ø �� 
͠          , 
^L 	;H 
j 	;H 
j 	n 
^L 	n 
^L 	;H          , 	 � 	;H 	h 	;H 	h 	�0 	 � 	�0 	 � 	;H          , +z� �\ +�� �\ +�� � +z� � +z� �\          , �� �� ְ �� ְ ߜ �� ߜ �� ��          , 	#� �h 	/� �h 	/� % 	#� % 	#� �h          , %T �( % �( % � %T � %T �(          , I� %�L U� %�L U� &3L I� &3L I� %�L          , T� % `� % `� &3L T� &3L T� %          , 
�  �� L  �� L X 
� X 
�  ��          ,  i� )� i� )� ø  ø  i�          , �� �� �� �� �� � �� � �� ��          , 4� � @p � @p C< 4� C< 4� �          , �H �� �  �� �  #I4 �H #I4 �H ��          , &�l �T &�$ �T &�$ � &�l � &�l �T          , '�P 0� '� 0� '� H� '�P H� '�P 0�          , 
h L 
s� L 
s� , 
h , 
h L          , ,�p �L ,�( �L ,�( V ,�p V ,�p �L          , � !x &� !x &� T@ � T@ � !x          , '��  ' '�d  ' '�d  Y� '��  Y� '��  '          , j� �� vp �� vp  Ơ j�  Ơ j� ��          , �� � �| � �| �� �� �� �� �          , � �4 �� �4 �� "� � "� � �4          , 	j( �L 	u� �L 	u� � 	j( � 	j( �L          , �X O � O � fd �X fd �X O          , � �� �H �� �H fd � fd � ��          , �� �d h �d h  ��  �� �d          , %7X �( %C �( %C �� %7X �� %7X �(          , 
͠  � 
�X  � 
�X � 
͠ � 
͠  �          , 
�x ( 
�0 ( 
�0 Z� 
�x Z� 
�x (          , "�( �4 "�� �4 "��   � "�(   � "�( �4          , *�h S� *�  S� *�  �t *�h �t *�h S�          , ,�p h ,�( h ,�( E0 ,�p E0 ,�p h          , (�� h (� h (� E0 (�� E0 (�� h          ,  zt $��  �, $��  �, %�  zt %�  zt $��          , .x| �� .�4 �� .�4 �� .x| �� .x| ��          , &5@  � &@�  � &@� �p &5@ �p &5@  �          , 0�( �� 1� �� 1� }d 0�( }d 0�( ��          , � � �d � �d �� � �� � �          , �� \ �� \ �� 	�X �� 	�X �� \          , )��  4� )�p  4� )�p �� )�� �� )��  4�          , &� 8T &�� 8T &�� k &� k &� 8T          ,  | ;� ,4 ;� ,4 ø  | ø  | ;�          , Q, 
`@ \� 
`@ \� _� Q, _� Q, 
`@          , *ڴ !�\ *�l !�\ *�l "($ *ڴ "($ *ڴ !�\          , /h %�L ;  %�L ;  &74 /h &74 /h %�L          ,  � 	f@ ,� 	f@ ,� �  � �  � 	f@          , $�H :� $�  :� $�  m� $�H m� $�H :�          , 0�( 7\ 1� 7\ 1� j$ 0�( j$ 0�( 7\          , )�H Đ )�  Đ )�  nX )�H nX )�H Đ          , *<�  � *H8  � *H8 �H *<� �H *<�  �          , 	�� 
� 
h 
� 
h �� 	�� �� 	�� 
�          , d� �4 p� �4 p� 	� d� 	� d� �4          , !� �� !�h �� !�h �� !� �� !� ��          , +�� �p +�8 �p +�8 f� +�� f� +�� �p          , ֈ �� �@ �� �@ �T ֈ �T ֈ ��          , �� eD �\ eD �\ �� �� �� �� eD          , � � @ � @ �� � �� � �          , -�l ~@ -�$ ~@ -�$ /H -�l /H -�l ~@          , � $ � $ � "($ � "($ � $          , 4L Đ @ Đ @ � 4L � 4L Đ          , $I 4P $T� 4P $T� �t $I �t $I 4P          , Rp  � ^(  � ^( X Rp X Rp  �          , *�( 0� *�� 0� *�� p� *�( p� *�( 0�          , 
D d� 
� d� 
� �� 
D �� 
D d�          , 'g� �� 's� �� 's� � 'g� � 'g� ��          , � �� l �� l ?� � ?� � ��          , %�� Y� %�� Y� %�� �� %�� �� %�� Y�          , Ah 	�� M  	�� M  �� Ah �� Ah 	��          , � 7� �� 7� �� � � � � 7�          , &�x �l '0 �l '0 �| &�x �| &�x �l          , а � �h � �h ?� а ?� а �          , �� "� �� "� �� #& �� #& �� "�          , �� "�D �h "�D �h #& �� #& �� "�D          , �� �� �x �� �x !� �� !� �� ��          , S� �\ _� �\ _� �| S� �| S� �\          , 0�( eD 1� eD 1� � 0�( � 0�( eD          , (X  �T (c� �T (c� �� (X  �� (X  �T          , '�  
� '�� 
� '�� =� '�  =� '�  
�          , $l8 
� $w� 
� $w� =� $l8 =� $l8 
�          , ?T !� K !� K #ݤ ?T #ݤ ?T !�          , �� d$ �| d$ �| �� �� �� �� d$          , �� �\ �T �\ �T +� �� +� �� �\          , $5� `< $A@ `< $A@ � $5� � $5� `<          , o� 	�P {P 	�P {P 	� o� 	� o� 	�P          , Ѩ 	�8 �` 	�8 �` I� Ѩ I� Ѩ 	�8          , &F� :l &R� :l &R� m4 &F� m4 &F� :l          , �t �8 �, �8 �, �| �t �| �t �8          , 	�� � 	�� � 	�� VT 	�� VT 	�� �          , ؀ !�T �8 !�T �8 !� ؀ !� ؀ !�T          , (!p  � (-(  � (-( �� (!p �� (!p  �          , "1� �� "=� �� "=� �| "1� �| "1� ��          , L �L W� �L W� � L � L �L          , 'm� [ 'yx [ 'yx m� 'm� m� 'm� [          , $X�  � $dh  � $dh @ $X� @ $X�  �          , ]� �( iP �( iP �� ]� �� ]� �(          ,  | S� ,4 S� ,4 �L  | �L  | S�          , �t �8 �, �8 �, )  �t )  �t �8          ,  6 �  A� �  A� �  6 �  6 �          , I8 4P T� 4P T� f� I8 f� I8 4P          , L� � X� � X� �� L� �� L� �          , /� �t ;h �t ;h �� /� �� /� �t          , 	� T@ 	�� T@ 	�� �| 	� �| 	� T@          , 	�l ;� 	�$ ;� 	�$ _� 	�l _� 	�l ;�          , (� 
( (�� 
( (�� �� (� �� (� 
(          , ' �T 2� �T 2� � ' � ' �T          , �\ H � H � ( �\ ( �\ H          , �� 	;H �h 	;H �h 	� �� 	� �� 	;H          , S� T@ _H T@ _H � S� � S� T@          , �X �� � �� � �� �X �� �X ��          , �T 3� � 3� � �� �T �� �T 3�          , :p 3� F( 3� F( f� :p f� :p 3�          , ~� �$ �� �$ �� !4  ~� !4  ~� �$          , "� 	?0 #� 	?0 #� � "� � "� 	?0          , (�< �� )� �� )�  (�<  (�< ��          , 	�� %�$ 	Ք %�$ 	Ք 'T 	�� 'T 	�� %�$          , �� 	� �� 	� �� <h �� <h �� 	�          , :�   FL   FL "�� :� "�� :�            ,   �  � iP  iP            , .$�  � .08  � .08 �� .$� �� .$�  �          , 6< � A� � A� 	� 6< 	� 6< �          , H< C\ S� C\ S� �| H< �| H< C\          , �8 v� �� v� �� �| �8 �| �8 v�          , )| ?t )%4 ?t )%4 � )| � )| ?t          , � $ +� $ +� �H � �H � $          , �  u0 ��  u0 �� ~� � ~� �  u0          , �  Z� �� Z� �� �t �  �t �  Z�          , $�  0� $�� 0� $�� p� $�  p� $�  0�          , 	!�  ' 	-�  ' 	-�  Y� 	!�  Y� 	!�  '          , �l Wx �$ Wx �$ �\ �l �\ �l Wx          , �8 &'� �� &'� �� &Z\ �8 &Z\ �8 &'�          , O�  �� [�  �� [� $-� O� $-� O�  ��          , �� ;� �| ;� �| �� �� �� �� ;�          , � ,� �� ,� �� q  � q  � ,�          , -|� �x -�@ �x -�@   -|�   -|� �x          , � z� �� z� ��   �   � z�          , �` H� � H� � % �` % �` H�          , I� � U8 � U8 � I� � I� �          , � =� � =� � �� � �� � =�          , S� � _� � _� Q S� Q S� �          , q� %�L }D %�L }D &Z\ q� &Z\ q� %�L          , )�� �� )� �� )� �� )�� �� )�� ��          , �<  �� ��  �� �� �  �< �  �<  ��          , �� #�� �� #�� �� &�l �� &�l �� #��          , �� /� �L /� �L nX �� nX �� /�          , ,�� � -d � -d �� ,�� �� ,�� �          , %�� �h %׀ �h %׀ ?� %�� ?� %�� �h          , h �   �   y4 h y4 h �          , �� �� ׬ �� ׬ !zP �� !zP �� ��          , 	/� "� 	;H "� 	;H #� 	/� #� 	/� "�          , :l , F$ , F$ !�� :l !�� :l ,          , � �� %� �� %� N@ � N@ � ��          , $հ %�  $�h %�  $�h 'T $հ 'T $հ %�           , -c$ �< -n� �< -n� �� -c$ �� -c$ �<          , ,.� �  ,:D �  ,:D �� ,.� �� ,.� �           , ,k � ,v� � ,v� p� ,k p� ,k �          , *� �� *d �� *d @( *� @( *� ��          , W� �� cp �� cp ۴ W� ۴ W� ��          , *�� :l +� :l +� �T *�� �T *�� :l          , $�@ L $�� L $�� �T $�@ �T $�@ L          , n0 :l y� :l y� m4 n0 m4 n0 :l          , '�X � '� � '� t� '�X t� '�X �          , $�h �4 $�  �4 $�  � $�h � $�h �4          , k� �� w� �� w� �@ k� �@ k� ��          , �\ �, � �, � �T �\ �T �\ �,          , ${� ȼ $�� ȼ $�� p� ${� p� ${� ȼ          , '� �l ''p �l ''p o� '� o� '� �l          , !�� �� !�d �� !�d ۴ !�� ۴ !�� ��          , - �D 8� �D 8� �d - �d - �D          , �H N� �  N� �  iL �H iL �H N�          , �\ Wx  Wx  t� �\ t� �\ Wx          , (P ٜ 4 ٜ 4 m4 (P m4 (P ٜ          , �` b� � b� � � �` � �` b�          , $�D �� $�� �� $�� �L $�D �L $�D ��          , Ŭ �P �d �P �d �4 Ŭ �4 Ŭ �P          , *[� \� *gx \� *gx �� *[� �� *[� \�          , )y0 � )�� � )�� pL )y0 pL )y0 �          , .� ;� ."� ;� ."� pL .� pL .� ;�          , .I� �< .UT �< .UT �� .I� �� .I� �<          , 	Ѭ � 	�d � 	�d   	Ѭ   	Ѭ �          , f� �� r� �� r� C< f� C< f� ��          , h $פ )  $פ )  %� h %� h $פ          , �� !�L �l !�L �l &�l �� &�l �� !�L          ,  � `  X `  X L(  � L(  � `          , z| J� �4 J� �4 s� z| s� z| J�          , � �� �8 �� �8 /D � /D � ��          , #H !�L #(  !�L #(  "($ #H "($ #H !�L          , $�p '< $�( '< $�( '%| $�p '%| $�p '<          , $݀ '� $�8 '� $�8 'L� $݀ 'L� $݀ '�          , �L 4 � 4 � 
�  �L 
�  �L 4          , &  �� &�  �� &� ! & ! &  ��          , �8 �  �� �  ��  � �8  � �8 �           , �� d� �l d� �l �p �� �p �� d�          , m �� x� �� x� �� m �� m ��          , �@ ( �� ( �� @ �@ @ �@ (          , �� �� �� �� �� ø �� ø �� ��          , Y� �� e� �� e� ?� Y� ?� Y� ��          , 'w�  � '�<  � '�< � 'w� � 'w�  �          , &�h  �� &�   �� &�  � &�h � &�h  ��          , )�T  � )�  � )� X )�T X )�T  �          , 9 7� D� 7� D� L( 9 L( 9 7�          , %�p �� %�( �� %�( �, %�p �, %�p ��          , .08 #�� .;� #�� .;� $� .08 $� .08 #��          , -�� #�� -�| #�� -�| $� -�� $� -�� #��          , \T � h � h �� \T �� \T �          , !l� z� !x\ z� !x\ nX !l� nX !l� z�          , #f� %�  #r8 %�  #r8 &d  #f� &d  #f� %�           , �0 O �� O �� �t �0 �t �0 O          , 
�@ � 
�� � 
�� jL 
�@ jL 
�@ �          , �P �L � �L �  Ơ �P  Ơ �P �L          , )�D � )�� � )�� �� )�D �� )�D �          , % �� 0� �� 0� �D % �D % ��          , � �� �� �� �� �D � �D � ��          , � �� �� �� �� F$ � F$ � ��          ,   � �  � � ��  ��   �          , )� 
�h 5h 
�h 5h � )� � )� 
�h          , $�X D $� D $� m4 $�X m4 $�X D          , v� �� �� �� �� 
�H v� 
�H v� ��          , � 	f@ �l 	f@ �l p� � p� � 	f@          , �P H � H � L( �P L( �P H          , �P 7� � 7� � j� �P j� �P 7�      >    , � $�� �� $�� �� $�< � $�< � $��      >    , �$ i� �  i� �  u� �$ u� �$ i�      >    , * �� W� �� W� �� * �� * ��      >    , P i� ,� i� ,� u� P u� P i�      >    , ?t �� x �� x �� ?t �� ?t ��      >    , �< $ y8 $ y8 "� �< "� �< $      >    , #� B� y8 B� y8 N@ #� N@ #� B�      >    ,  � 	f@  � 	f@  � 	q�  � 	q�  � 	f@      >    , | ;� �� ;� �� GH | GH | ;�      >    , �� $�� �h $�� �h $�d �� $�d �� $��      >    ,  � �8 �L �8 �L �  � �  � �8      >    , -A� �� -p� �� -p� �� -A� �� -A� ��      >    , m� �� L �� L �� m� �� m� ��      >    , )�H b� *!( b� *!( nX )�H nX )�H b�      >    , )�� � *� � *� �� )�� �� )�� �      >    , �P �L #� �L #� � �P � �P �L      >    , '�� �� (H� �� (H� �D '�� �D '�� ��      >    , '�� �| )>� �| )>� �4 '�� �4 '�� �|      >    , %� �T &`8 �T &`8 � %� � %� �T      >    , �D &'� � &'� � &3L �D &3L �D &'�      >    , &1X 0� '� 0� '� <d &1X <d &1X 0�      >    , %bP �@ %Ә �@ %Ә �� %bP �� %bP �@      >    , &��  � ' `  � ' `  d &��  d &��  �      >    , #T   $l   $l � #T � #T        >    , $� ', %�� ', %�� 2� $� 2� $� ',      >    , q  ٜ �� ٜ �� �T q  �T q  ٜ      >    , �4 't  't  3, �4 3, �4 't      >    , +]� Z� -p� Z� -p� f� +]� f� +]� Z�      >    , -A� �� -p� �� -p� Ӝ -A� Ӝ -A� ��      >    , .UT � .�4 � .�4 �� .UT �� .UT �      >    , �@ !�L � !�L � !� �@ !� �@ !�L      >    , x� �� $G �� $G �� x� �� x� ��      >    , $?L �� 1� �� 1� �� $?L �� $?L ��      >    , *@ ( ,�� ( ,�� � *@ � *@ (      >    , (�p �� )�� �� )�� �� (�p �� (�p ��      >    , '�� = (�( = (�( H� '�� H� '�� =      >    , �\ �� �� �� �� �\ �\ �\ �\ ��      >    , !A� �4 "� �4 "� �� !A� �� !A� �4      >    , %�� � &�� � &�� �� %�� �� %�� �      >    , �X 0�  � 0�  � <d �X <d �X 0�      >    , �� #�� � #�� � #� �� #� �� #��      >    , 
}� �8 � �8 � � 
}� � 
}� �8      >    , p( 
�� 	�8 
�� 	�8 \ p( \ p( 
��      >    , ��  �� �(  �� �(  �8 ��  �8 ��  ��      >    , �P d� � d� � pl �P pl �P d�      >    , *�h �� -d �� -d �t *�h �t *�h ��      >    ,  zt qh !� qh !� }   zt }   zt qh      >    , �P $Ӽ �� $Ӽ �� $�t �P $�t �P $Ӽ      >    , �, �4 L �4 L �� �, �� �, �4      >    , �� !�\ �� !�\ �� " �� " �� !�\      >    , O�  �� ��  �� ��  Ơ O�  Ơ O�  ��      >    , �� μ #�  μ #�  �t �� �t �� μ      >    , "�� �� $)� �� $)� �� "�� �� "�� ��      >    , $"  �� %N� �� %N� �� $"  �� $"  ��      >    , #�, μ .[0 μ .[0 �t #�, �t #�, μ      >    , )�X i, *Y� i, *Y� t� )�X t� )�X i,      >    , *.� v� *_� v� *_� �� *.� �� *.� v�      >    , �� d$ �| d$ �| o� �� o� �� d$      >    , q�  ' ��  ' ��  2� q�  2� q�  '      >    , ��  ' 	-�  ' 	-�  2� ��  2� ��  '      >    , i0  ' ��  ' ��  2� i0  2� i0  '      >    , )8� 0� *�� 0� *�� <d )8� <d )8� 0�      >    , �` #� (� #� (� /D �` /D �` #�      >    , �� �� �� �� �� � �� � �� ��      >    , �  � �� � �� �� �  �� �  �      >    , 	�  �4 	�  �4 	�  �� 	�  �� 	�  �4      >    , 	3x ;� 	Ӡ ;� 	Ӡ GH 	3x GH 	3x ;�      >    , :l , "f� , "f�  � :l  � :l ,      >    , a< %�\ �  %�\ �  %� a< %� a< %�\      >    , +M� #� +�� #� +�� /D +M� /D +M� #�      >    , '�� `< +Y� `< +Y� k� '�� k� '�� `<      >    , μ d� �D d� �D p� μ p� μ d�      >    , E� �� t� �� t� �� E� �� E� ��      >    , ?� �T �d �T �d � ?� � ?� �T      >    , 4P :l p� :l p� F$ 4P F$ 4P :l      >    , �4 �� � �� � ڔ �4 ڔ �4 ��      >    , (-( �@ (�( �@ (�( �� (-( �� (-( �@      >    , �� ٜ �� ٜ �� �T �� �T �� ٜ      >    , 0 �, �� �, �� �� 0 �� 0 �,      >    , *� ȼ ,� ȼ ,� �t *� �t *� ȼ      >    , *� �� +�� �� +�� �� *� �� *� ��      >    , �� �� �d �� �d �\ �� �\ �� ��      >    , ݬ m|   m|   y4 ݬ y4 ݬ m|      >    , �h �� *� �� *� �D �h �D �h ��      >    , "� `<  �@ `<  �@ k� "� k� "� `<      >    , �� �4 7� �4 7� �� �� �� �� �4      >    , �� "� ߜ "� ߜ "�� �� "�� �� "�      >    , z| J� 9� J� 9� VT z| VT z| J�      >    , '� C V� C V� N� '� N� '� C      >    , � �� p �� p �T � �T � ��      >    , *�( d� *�` d� *�` p� *�( p� *�( d�      >    , �  �� �  �� �  �8 �  �8 �  ��      >    , "~ �4 "�� �4 "�� �� "~ �� "~ �4      >    , r< d� �� d� �� pl r< pl r< d�      >    , �� �| �� �| �� �4 �� �4 �� �|      >    , ,$� �� -�� �� -�� �� ,$� �� ,$� ��      >    , �� ', � ', � 2� �� 2� �� ',      >    , !4  �8 !�@ �8 !�@ � !4  � !4  �8      >    ,  �� �8 !5� �8 !5� �  �� �  �� �8      >    , I� �� h� �� h� �T I� �T I� ��      >    , � ʬ �� ʬ �� �d � �d � ʬ      >    ,  8� :l t� :l t� F$  8� F$  8� :l      >    , 	#� � 	s� � 	s� < 	#� < 	#� �      >    , 	H� 8T �� 8T �� D 	H� D 	H� 8T      >    , y� d� �� d� �� p� y� p� y� d�      >    ,  �  �  �  �  �  �X  �  �X  �  �      >    , #(  d� #V� d� #V� pl #(  pl #(  d�      >    , �� �| *� �| *� �4 �� �4 �� �|      >    , � �� M� �� M� �t � �t � ��      >    , �� [ f� [ f� f� �� f� �� [      >    , ��  � �  � �  �H ��  �H ��  �      >    , )+ 	�x +� 	�x +� 	�0 )+ 	�0 )+ 	�x      >    , %�� 	�x )- 	�x )- 	�0 %�� 	�0 %�� 	�x      >    , P $�� 	� $�� 	� $�L P $�L P $��      >    , 'ˀ 	� (B� 	� (B� x 'ˀ x 'ˀ 	�      >    , (%X �� )� �� )� �L (%X �L (%X ��      >    , � � p  � p  �� � �� � �      >    , ',  d ��  d ��  ',  ',  d      >    , Qt � &= � &= < Qt < Qt �      >    , !� 4 "?� 4 "?� ?� !� ?� !� 4      >    , �� �� �h �� �h �� �� �� �� ��      >    , �t !� W� !� W� !�� �t !�� �t !�      >    , *ܨ �� ,�8 �� ,�8 �L *ܨ �L *ܨ ��      >    , *�@ #� *�T #� *�T /D *�@ /D *�@ #�      >    , #H Ll %�� Ll %�� X$ #H X$ #H Ll      >    , "�� 	f@ #t, 	f@ #t, 	q� "�� 	q� "�� 	f@      >    , #r8 	f@ $�� 	f@ $�� 	q� #r8 	q� #r8 	f@      >    ,  d �� � �� � �D  d �D  d ��      >    , )�X � )�  � )�  � )�X � )�X �      >    , %�� �� 'i� �� 'i� �� %�� �� %�� ��      >    , (P 	f@  	f@  	q� (P 	q� (P 	f@      >    , 1� 4 �� 4 �� ?� 1� ?� 1� 4      >    , $� �0 $�� �0 $�� �� $� �� $� �0      >    , ,k d� ,�  d� ,�  p� ,k p� ,k d�      >    , 4� 
d( x� 
d( x� 
o� 4� 
o� 4� 
d(      >    , 4� �� ؤ �� ؤ ٠ 4� ٠ 4� ��      >    , &l �X (� �X (� � &l � &l �X      >    , l�   1�   1� � l� � l�        >    , W0 "^� Ex "^� Ex "j� W0 "j� W0 "^�      >    , �l !�\ "P !�\ "P " �l " �l !�\      >    , +q >4 +�, >4 +�, I� +q I� +q >4      >    , +�t eD -|� eD -|� p� +�t p� +�t eD      >    , �� `< � `< � k� �� k� �� `<      >    , �h  ' f�  ' f�  2� �h  2� �h  '      >    , �h � x� � x� �� �h �� �h �      >    , R( ;� � ;� � GH R( GH R( ;�      >    , ^ ;� T ;� T GH ^ GH ^ ;�      >    , %�  � �L  � �L  �H %�  �H %�  �      >    , �l Wx �L Wx �L c0 �l c0 �l Wx      >    , �� �� �� �� �� �� �� �� �� ��      >    , ?P �, �� �, �� �� ?P �� ?P �,      >    , "M@ x *<� x *<� '0 "M@ '0 "M@ x      >    , (�� eD )�( eD )�( p� (�� p� (�� eD      >    , � ~@ ]L ~@ ]L �� � �� � ~@      >    , �|  �� .(  �� .(  �8 �|  �8 �|  ��      >    , ^H :l �L :l �L F$ ^H F$ ^H :l      >    , _$ !�< SH !�< SH !�� _$ !�� _$ !�<      >    , ,� !�< a !�< a !�� ,� !�� ,� !�<      >    , %Ѥ =� '5 =� '5 I� %Ѥ I� %Ѥ =�      >    , � d� � d� � p� � p� � d�      >    , �( ~@ 	� ~@ 	� �� �( �� �( ~@      >    , �� 4 3 4 3 ?� �� ?� �� 4      >    , x` �� �� �� �� �L x` �L x` ��      >    , � �� ~` �� ~` �D � �D � ��      >    , \ �� �  �� �  �| \ �| \ ��      >    , f� �� ;� �� ;� �t f� �t f� ��      >    , H� !�L Jx !�L Jx !� H� !� H� !�L      >    , -� �8 �� �8 �� � -� � -� �8      >    , �� S� � S� � _� �� _� �� S�      >    , *B\ � ,t� � ,t�  8 *B\  8 *B\ �      >    , �@ #�� �  #�� �  #� �@ #� �@ #��      >    , e� ";� qd ";� qd "Gd e� "Gd e� ";�      >    , e� !`�  � !`�  � !l� e� !l� e� !`�      >    , �� \ �P \ �P  ��  �� \      >    , �� �� �  �� �  ڔ �� ڔ �� ��      >    , �P $jD T $jD T $u� �P $u� �P $jD      >    , � �� �8 �� �8 �D � �D � ��      >    , ., �X S$ �X S$ � ., � ., �X      >    , �L ;� � ;� � GH �L GH �L ;�      >    , g� i� �� i� �� u� g� u� g� i�      >    , %� |� &@� |� &@� �p %� �p %� |�      >    , 	�X :l XL :l XL F$ 	�X F$ 	�X :l      >    , !�  
d( !�� 
d( !�� 
o� !�  
o� !�  
d(      >    ,  �0 ;� !� ;� !� GH  �0 GH  �0 ;�      >    , -p �� -I� �� -I� �t -p �t -p ��      >    , ( :l �8 :l �8 F$ ( F$ ( :l      >    , �� !=� 4 !=� 4 !I| �� !I| �� !=�      >    , 4 6< |� 6< |� A� 4 A� 4 6<      >    , r� :l <  :l <  F$ r� F$ r� :l      >    , 
1` �� }h �� }h �D 
1` �D 
1` ��      >    , %� �0 	/� �0 	/� �� %� �� %� �0      >    , % � �� %�� �� %�� �D % � �D % � ��      >    , #۰ 4 $^� 4 $^� ?� #۰ ?� #۰ 4      >    , �| �8 �P �8 �P � �| � �| �8      >    , v� �8 �� �8 �� � v� � v� �8      >    , %� �@ &%� �@ &%� �� %� �� %� �@      >    , �l ȼ !S@ ȼ !S@ �t �l �t �l ȼ      >    , |$ 	f@ �| 	f@ �| 	q� |$ 	q� |$ 	f@      >    , �� �| �d �| �d �4 �� �4 �� �|      >    , � �P � �P � � � � � �P      >    , �� 4P '� 4P '� @ �� @ �� 4P      >    , 
�< �| �T �| �T �4 
�< �4 
�< �|      >    , &�< � ()@ � ()@ �p &�< �p &�< �      >    ,  =� �T !I| �T !I| �  =� �  =� �T      >    , �  �h �( �h �( �  �  �  �  �h      >    , e� 	 q@ 	 q@ 	'� e� 	'� e� 	      >    , 1  � 	�  � 	�  �H 1  �H 1  �      >    , #� � 	� � 	� �� #� �� #� �      >    , -&� �� -� �� -� � -&� � -&� ��      >    , �� !� �� !� �� !�� �� !�� �� !�      >    , 	1� :l 	�L :l 	�L F$ 	1� F$ 	1� :l      >    , �H #=|  � #=|  � #I4 �H #I4 �H #=|      >    , "� %�\ "�T %�\ "�T %� "� %� "� %�\      >    , VT   o�   o� � VT � VT        >    , %�h �x &� �x &� �0 %�h �0 %�h �x      >    , �< �| 2� �| 2� �4 �< �4 �< �|      >    , Y� �� &� �� &� �p Y� �p Y� ��      >    , �� � 1� � 1� %\ �� %\ �� �      >    , `   U8   U8 � ` � `        >    , ,�� �T -�t �T -�t � ,�� � ,�� �T      >    , b� c� �p c� �p oL b� oL b� c�      >    , +"� �T ,� �T ,� � +"� � +"� �T      >    , Z�  �� t  �� t  �8 Z�  �8 Z�  ��      >    ,  | �� W, �� W, �L  | �L  | ��      >    , �h }� �H }� �H �� �h �� �h }�      >    , �| !� �  !� �  !�� �| !�� �| !�      >    , )�� :l *�� :l *�� F$ )�� F$ )�� :l      >    , U| ^�  � ^�  � jL U| jL U| ^�      >    , � �P  � �P  � 
 � 
 � �P      >    , B� �� � �� � �� B� �� B� ��      >    , 
� ٜ �H ٜ �H �T 
� �T 
� ٜ      >    , T� �� �� �� �� �@ T� �@ T� ��      >    , \� �� X� �� X� < \� < \� ��      >    , p( &l � &l � &$ p( &$ p( &l      >    , N< x� �� x� �� �\ N< �\ N< x�      >    ,   Ll #< Ll #< X$   X$   Ll      >    , �� � �� � �� �� �� �� �� �      >    , 	�� %�$ 	Ք %�$ 	Ք %�� 	�� %�� 	�� %�$      >    , '�X 	f@ (X  	f@ (X  	q� '�X 	q� '�X 	f@      >    , (PP � -0\ � -0\ �� (PP �� (PP �      >    , %�� 4 &� 4 &� ?� %�� ?� %�� 4      >    , � ?t %� ?t %� K, � K, � ?t      >    , �L H T H T )  �L )  �L H      >    , � �  �  �p � �p � �      >    , $l  �� %�  �� %�  �8 $l  �8 $l  ��      >    , � ,�  �� ,�  �� 8� � 8� � ,�      >    , L( 4 � 4 � ?� L( ?� L( 4      >    , X 4 N 4 N ?� X ?� X 4      >    , �( "� 
s� "� 
s� "�� �( "�� �( "�      >    , %�( �� (�$ �� (�$ �� %�( �� %�( ��      >    , %�\ �8 &�  �8 &�  � %�\ � %�\ �8      >    , %�0 eD &� eD &� p� %�0 p� %�0 eD      >    , %�� � &ˤ � &ˤ  8 %��  8 %�� �      >    , #
� 	�x %f8 	�x %f8 	�0 #
� 	�0 #
� 	�x      >    , )	� %�\ *FD %�\ *FD %� )	� %� )	� %�\      >    , ʌ �4   �4   �� ʌ �� ʌ �4      >    , E0 !n� ׬ !n� ׬ !zP E0 !zP E0 !n�      >    , (� >4 �� >4 �� I� (� I� (� >4      >    , U8 �� � �� � �� U8 �� U8 ��      >    , � Đ � Đ � �H � �H � Đ      >    , �� Đ � Đ � �H �� �H �� Đ      >    , 2� d� � d� � p� 2� p� 2� d�      >    , )�� �  *(� �  *(� �� )�� �� )�� �       >    , #H �� #�� �� #�� �� #H �� #H ��      >    , �t  #(   #(   � �t  � �t       >    , � !�\ - !�\ - " � " � !�\      >    , �� :l a� :l a� F$ �� F$ �� :l      >    , )�D >4 *d >4 *d I� )�D I� )�D >4      >    , �� �T �p �T �p � �� � �� �T      >    ,  � c� I� c� I� oP  � oP  � c�      >    , 
� $  � $  � $+� 
� $+� 
� $       >    , � 	?0 �| 	?0 �| 	J� � 	J� � 	?0      >    , U| ~@ #f� ~@ #f� �� U| �� U| ~@      >    , 	\| � 
� � 
� �� 	\| �� 	\| �      >    , �0 � 	^p � 	^p �� �0 �� �0 �      >    , $�( Y� &�� Y� &�� eH $�( eH $�( Y�      >    , �� �| �� �| �� �4 �� �4 �� �|      >    ,  0< ��  �� ��  �� ��  0< ��  0< ��      >    , *�X U` *�x U` *�x a *�X a *�X U`      >    , !� #�� #�@ #�� #�@ $� !� $� !� #��      >    , *� �8 +�  �8 +�  � *� � *� �8      >    , WP 	f@ �l 	f@ �l 	q� WP 	q� WP 	f@      >    , #�h :l $�8 :l $�8 F$ #�h F$ #�h :l      >    , �� :l  p� :l  p� F$ �� F$ �� :l      >    , 	H� !$` 	w� !$` 	w� !0 	H� !0 	H� !$`      >    , �� �� 	 �� 	 �T �� �T �� ��      >    , '� �l ,r� �l ,r� �$ '� �$ '� �l      >    , &+| �D &�� �D &�� �� &+| �� &+| �D      >    , �� $ � �x $ � �x $� �� $� �� $ �      >    , *Q� >4 +.� >4 +.� I� *Q� I� *Q� >4      >    , b� 	� dH 	� dH X b� X b� 	�      >    , �d �h �$ �h �$ �  �d �  �d �h      >    , m #�� � #�� � $� m $� m #��      >    , yX #�� �( #�� �( #� yX #� yX #��      >    , R� %�L s� %�L s� %� R� %� R� %�L      >    , �� �T �� �T �� � �� � �� �T      >    , �� �T �@ �T �@ � �� � �� �T      >    , -�� �� 1� �� 1� �� -�� �� -�� ��      >    , +�4 �� ,&� �� ,&� �� +�4 �� +�4 ��      >    , �( �T �� �T �� � �( � �( �T      >    , �� �T �� �T �� � �� � �� �T      >    , "�� d� "�p d� "�p pl "�� pl "�� d�      >    , %#� b� &@� b� &@� nX %#� nX %#� b�      >    , &5@ ;� 'u� ;� 'u� GH &5@ GH &5@ ;�      >    , �� [ � [ � f� �� f� �� [      >    , �� O� e� O� e� [< �� [< �� O�      >    , � ;� 5� ;� 5� GH � GH � ;�      >    , 2| �� S� �� S� �D 2| �D 2| ��      >    , � !�\ K� !�\ K� " � " � !�\      >    , x< �$ �  �$ �  � x< � x< �$      >    , �l � ,6\ � ,6\ %� �l %� �l �      >    , #� �T $0 �T $0 � #� � #� �T      >    , *� ʬ &� ʬ &� �d *� �d *� ʬ      >    , �� �� w@ �� w@ < �� < �� ��      >    , 
!� �� 8 �� 8 �� 
!� �� 
!� ��      >    , %�� m| )B� m| )B� y4 %�� y4 %�� m|      >    , ,| �� ,6\ �� ,6\ �| ,| �| ,| ��      >    , y4 &�� |� &�� |� 'T y4 'T y4 &��      >    , ,� 4 ,�� 4 ,�� ?� ,� ?� ,� 4      >    , �� !�L �L !�L �L !� �� !� �� !�L      >    , � !� ހ !� ހ !�� � !�� � !�      >    , , "b� �$ "b� �$ "nt , "nt , "b�      >    , ,p� �| .WH �| .WH �4 ,p� �4 ,p� �|      >    , )$ d� �� d� �� pl )$ pl )$ d�      >    , z 
A  
� 
A  
� 
L� z 
L� z 
A       >    , �� :l �\ :l �\ F$ �� F$ �� :l      >    , �< !$` � !$` � !0 �< !0 �< !$`      >    , � a|   a|   m4 � m4 � a|      >    , �� a| � a| � m4 �� m4 �� a|      >    , !  ި O�  ި O�  �` !  �` !  ި      >    , "�� �� '� �� '� �t "�� �t "�� ��      >    , | �� � �� � �x | �x | ��      >    , �P %` �, %` �, 1 �P 1 �P %`      >    , !�� i� #� i� #� u� !�� u� !�� i�      >    , 9� �l �� �l �� $ 9� $ 9� �l      >    , � ', O� ', O� 2� � 2� � ',      >    , $� � %#� � %#� �< $� �< $� �      >    , $�  
� &!� 
� &!� 
)� $�  
)� $�  
�      >    , #+� a\ #z a\ #z m #+� m #+� a\      >    , #nP �� #�� �� #�� �� #nP �� #nP ��      >    , �� �� �  �� �  �� �� �� �� ��      >    , �, 	�  h 	�  h X �, X �, 	�      >    , I\   ��   �� � I\ � I\        >    , #b� �� $0 �� $0 �D #b� �D #b� ��      >    , �� #�� A  #�� A  $� �� $� �� #��      >    , � ', ?� ', ?� 2� � 2� � ',      >    , �| c�  O| c�  O| oL �| oL �| c�      >    , � �, 6� �, 6� �� � �� � �,      >    , ${� 
ш %׀ 
ш %׀ 
�@ ${� 
�@ ${� 
ш      >    , �� #�� �H #�� �H $� �� $� �� #��      >    , i0 	f@ Q� 	f@ Q� 	q� i0 	q� i0 	f@      >    , 
P� �� 
� �� 
� �� 
P� �� 
P� ��      >    , "�� � #f� � #f� �p "�� �p "�� �      >    , � :l �� :l �� F$ � F$ � :l      >    , )h �8 � �8 � � )h � )h �8      >    , �� \ ݨ \ ݨ  ��  �� \      >    , � �  A� �  A� �� � �� � �      >    , i(  � ��  � ��  �H i(  �H i(  �      >    , ڔ � � � � �� ڔ �� ڔ �      >    , e� � �� � �� (� e� (� e� �      >    , *�� z� *ڴ z� *ڴ �� *�� �� *�� z�      >    , +� �� ,|� �� ,|� �D +� �D +� ��      >    ,  6 N@ "� N@ "� Y�  6 Y�  6 N@      >    , � \ � \ �  �  � \      >    , � =�  =�  I� � I� � =�      >    , �< Z� � Z� � fd �< fd �< Z�      >    , �� 	�� �\ 	�� �\ 	�8 �� 	�8 �� 	��      >    , �� $ �� $ �� "� �� "� �� $      >    , *�@ ~@ - ~@ - �� *�@ �� *�@ ~@      >    , � !�L (� !�L (� !� � !� � !�L      >    , �  � ܈ � ܈ �� �  �� �  �      >    , .p =� �@ =� �@ I� .p I� .p =�      >    , Ќ >4 �h >4 �h I� Ќ I� Ќ >4      >    , ]� � m8 � m8 �� ]� �� ]� �      >    , X� L �h L �h ( X� ( X� L      >    , %!� �  'q� �  'q� ø %!� ø %!� �       >    , D 4 �� 4 �� ?� D ?� D 4      >    , �X ��   ��   �� �X �� �X ��      >    , �� �� �( �� �( �� �� �� �� ��      >    , zT #l �4 #l �4 #"$ zT #"$ zT #l      >    , � "�D �h "�D �h "�� � "�� � "�D      >    , �� U| "�\ U| "�\ a4 �� a4 �� U|      >    , � %�\ hT %�\ hT %� � %� � %�\      >    , �| � K � K �� �| �� �| �      >    , ,2t �� 1� �� 1� �� ,2t �� ,2t ��      >    ,  �� �h �� �h ��  ��  ��      >    , l 	� � 	� � X l X l 	�      >    , �H #�  �� #�  �� /D �H /D �H #�      >    , �8 !x &� !x &� -0 �8 -0 �8 !x      >    , @ �8 Z� �8 Z� � @ � @ �8      >    , !�h  d "�@  d "�@  !�h  !�h  d      >    , � $f\ �� $f\ �� $r � $r � $f\      >    , �T $C4 p $C4 p $N� �T $N� �T $C4      >    , _D 	?0 �� 	?0 �� 	J� _D 	J� _D 	?0      >    , � �� #�� �� #�� �| � �| � ��      >    , %�l � '{l � '{l �� %�l �� %�l �      >    , .� ( �� ( �� � .� � .� (      >    , #?p 4P $�d 4P $�d @ #?p @ #?p 4P      >    , /  !Kp ̤ !Kp ̤ !W( /  !W( /  !Kp      >    , �� �� �� �� �� �l �� �l �� ��      >    , .� S� !�( S� !�( _� .� _� .� S�      >    , %�� �P &R� �P &R� � %�� � %�� �P      >    , а � 9� � 9� � а � а �      >    , #b� ʬ #�0 ʬ #�0 �d #b� �d #b� ʬ      >    ,  	f@ C� 	f@ C� 	q�  	q�  	f@      >    ,  � _D � _D �p  �p  �      >    , S� � V� � V� �� S� �� S� �      >    , #�� �� %s� �� %s� �� #�� �� #�� ��      >    , zx 
�� =� 
�� =� 
�H zx 
�H zx 
��      >    , � �8 �� �8 �� � � � � �8      >    , |$ 7� �� 7� �� C< |$ C< |$ 7�      >    , 
� 28 9 28 9 =� 
� =� 
� 28      >    , �P 28 L 28 L =� �P =� �P 28      >    , � >4 d� >4 d� I� � I� � >4      >    , P� ;� �L ;� �L GH P� GH P� ;�      >    , K� ;� 6  ;� 6  GH K� GH K� ;�      >    , h %�\ 8 %�\ 8 %� h %� h %�\      >    , 	� L 	�� L 	�� ( 	� ( 	� L      >    , #� 
`@ �� 
`@ �� 
k� #� 
k� #� 
`@      >    , (�D h (� h (�   (�D   (�D h      >    , =� 	f@ � 	f@ � 	q� =� 	q� =� 	f@      >    , �� f< qh f< qh q� �� q� �� f<      >    , � �� �h �� �h �D � �D � ��      >    , \� "?� +\ "?� +\ "KL \� "KL \� "?�      >    , #\� |� $l8 |� $l8 �D #\� �D #\� |�      >    , Z� 	�x �� 	�x �� 	�0 Z� 	�0 Z� 	�x      >    , &�� \ (� \ (�  &��  &�� \      >    , &�� t &�� t &�� , &�� , &�� t      >    , ֈ  d h  d h  ֈ  ֈ  d      >    , s\ x �L x �L '0 s\ '0 s\ x      >    , b� � ", � ", $d b� $d b� �      >    , Fl d� �h d� �h pl Fl pl Fl d�      >    , 
h t 
�� t 
�� , 
h , 
h t      >    , Ŭ �P �� �P ��  Ŭ  Ŭ �P      >    , -A� �� .	( �� .	( �� -A� �� -A� ��      >    , Լ d� _h d� _h p� Լ p� Լ d�      >    , �4 ٜ �� ٜ �� �T �4 �T �4 ٜ      >    , �4 C �p C �p N� �4 N� �4 C      >    , 'T\ @ (�$ @ (�$ $� 'T\ $� 'T\ @      >    ,  �P eD !vh eD !vh p�  �P p�  �P eD      >    , #?p !�L $%� !�L $%� !� #?p !� #?p !�L      >    , ;D 	f@ �� 	f@ �� 	q� ;D 	q� ;D 	f@      >    , y 84 �� 84 �� C� y C� y 84      >    , /� � hT � hT �� /� �� /� �      >    , ,� �h b� �h b� �  ,� �  ,� �h      >    , �� � �� � �� � �� � �� �      >    , 2� � �� � �� �X 2� �X 2� �      >    , �� �� �` �� �` �� �� �� �� ��      >    , %� !�\ �� !�\ �� " %� " %� !�\      >    , ,� d� ܌ d� ܌ p� ,� p� ,� d�      >    , >0 d� g d� g p� >0 p� >0 d�      >    , k� ո �l ո �l �p k� �p k� ո      >    , D � ` � ` !t D !t D �      >    , !� ;� �� ;� �� G� !� G� !� ;�      >    , ְ ʬ � ʬ � �d ְ �d ְ ʬ      >    , �P #�� �` #�� �` $� �P $� �P #��      >    , p 	�� O` 	�� O` 	�` p 	�` p 	��      >    , � 
�` @ 
�` @ 
� � 
� � 
�`      >    , �� "b� �� "b� �� "nt �� "nt �� "b�      >    , � d� !P d� !P p� � p� � d�      >    , ! �� "5� �� "5� �� ! �� ! ��      >    , )Fh �T )�� �T )�� � )Fh � )Fh �T      >    , ƀ $f\ � $f\ � $r ƀ $r ƀ $f\      >    , ld a| `� a| `� m4 ld m4 ld a|      >    , %H� �( *@h �( *@h �� %H� �� %H� �(      >    , &� �� &ό �� &ό �� &� �� &� ��      >    , \T � H� � H� �� \T �� \T �      >    , �� $#� �d $#� �d $/� �� $/� �� $#�      >    , �( �� x� �� x� � �( � �( ��      >    , � 	�x #  	�x #  	�0 � 	�0 � 	�x      >    , � �� ^� �� ^� �� � �� � ��      >    , �,  �� �(  �� �(  �8 �,  �8 �,  ��      >    , y�  � L  � L  �H y�  �H y�  �      >    , ��  � {�  � {�  �H ��  �H ��  �      >    , +�� �  ,r� �  ,r� ø +�� ø +�� �       >    , +�t ٜ -�� ٜ -�� �T +�t �T +�t ٜ      >    , �� ;� [� ;� [� GH �� GH �� ;�      >    , ڼ ;� �� ;� �� GH ڼ GH ڼ ;�      >    , 	�x 	 J� 	 J� 	'� 	�x 	'� 	�x 	      >    , ~� "l � "l � "($ ~� "($ ~� "l      >    , �p � i, � i, � �p � �p �      >    , � "� �� "� �� "$< � "$< � "�      >    , +4� �� +gT �� +gT �T +4� �T +4� ��      >    , r� � � � � �� r� �� r� �      >    , H �� � �� � �| H �| H ��      >    , :p Z� �� Z� �� f� :p f� :p Z�      >    , �0 �  }@ �  }@ �� �0 �� �0 �       >    , !� i� �h i� �h u� !� u� !� i�      >    , �� !$` R� !$` R� !0 �� !0 �� !$`      >    , [< >X 3� >X 3� J [< J [< >X      >    , �X a| �8 a| �8 m4 �X m4 �X a|      >    , �0 � �H � �H �� �0 �� �0 �      >    , '�X �� (X  �� (X  �T '�X �T '�X ��      >    , � �� � �� � �� � �� � ��      >    , pL !Kp �� !Kp �� !W( pL !W( pL !Kp      >    , 4P $�l �\ $�l �\ $�$ 4P $�$ 4P $�l      >    , | � �� � �� �� | �� | �      >    , o, %�L U� %�L U� %� o, %� o, %�L      >    , �( &'� >0 &'� >0 &3L �( &3L �( &'�      >    , �0 &'� �  &'� �  &3L �0 &3L �0 &'�      >    , ,o  4� -| 4� -| @L ,o  @L ,o  4�      >    , P| � �( � �( � P| � P| �      >    , �( �( *d �( *d �� �( �� �( �(      >    , 3t n� bT n� bT zx 3t zx 3t n�      >    , V� �4 #� �4 #� �� V� �� V� �4      >    , �� =� �$ =� �$ I� �� I� �� =�      >    , �� !�<  l� !�<  l� !�� �� !�� �� !�<      >    , Xl H �L H �L )  Xl )  Xl H      >    , Mh ;� `� ;� `� GH Mh GH Mh ;�      >    , #�� �� %�$ �� %�$ �| #�� �| #�� ��      >    , �0 !�< � !�< � !�� �0 !�� �0 !�<      >    , 	, >4 
90 >4 
90 I� 	, I� 	, >4      >    , 
^L  d ��  d ��  
^L  
^L  d      >    , �p �| �T �| �T �4 �p �4 �p �|      >    , �  �� � �� � �| �  �| �  ��      >    , "( d� p d� p p� "( p� "( d�      >    , 0� �( iP �( iP �� 0� �� 0� �(      >    , & H � H � )  & )  & H      >    , ( a| 4 a| 4 m4 ( m4 ( a|      >    , X |� )h |� )h �D X �D X |�      >    , ~�  d ��  d ��  ~�  ~�  d      >    , 	��   
?   
? � 	�� � 	��        >    , %�0 !�< &͘ !�< &͘ !�� %�0 !�� %�0 !�<      >    , �� >4 �� >4 �� I� �� I� �� >4      >    , �| � : � : �� �| �� �| �      >    , "� �� #CX �� #CX �� "� �� "� ��      >    , l� #�� !�� #�� !�� $� l� $� l� #��      >    , �h  � `�  � `�  �H �h  �H �h  �      >    , %^h �� &F� �� &F� �T %^h �T %^h ��      >    , � !�< �� !�< �� !�� � !�� � !�<      >    , P &l �� &l �� &$ P &$ P &l      >    , Լ H Yh H Yh )  Լ )  Լ H      >    , �� �  rd �  rd ø �� ø �� �       >    , Rp � }h � }h �� Rp �� Rp �      >    , �� � �l � �l < �� < �� �      >    , �� $ �� $ �� "� �� "� �� $      >    , �D ?x ^$ ?x ^$ K0 �D K0 �D ?x      >    , l Z� �� Z� �� fd l fd l Z�      >    , 4� Đ �@ Đ �@ �H 4� �H 4� Đ      >    , ]� �8 �d �8 �d � ]� � ]� �8      >    , 	�� =� 
A  =� 
A  I� 	�� I� 	�� =�      >    , }� �� �� �� �� �D }� �D }� ��      >    , D ]� 5$ ]� 5$ iL D iL D ]�      >    , {P S� a� S� a� _� {P _� {P S�      >    , �� d� �p d� �p p� �� p� �� d�      >    , �� ^� X ^� X j� �� j� �� ^�      >    , #�� `< $A@ `< $A@ k� #�� k� #�� `<      >    , %��  d ':�  d ':�  %��  %��  d      >    , (��  � )�  � )�  �H (��  �H (��  �      >    , %�P  �� '�@  �� '�@  � %�P  � %�P  ��      >    , �` ` 	/� ` 	/� % �` % �` `      >    , 	#� �h 
�� �h 
�� �  	#� �  	#� �h      >    , $hP �� %�� �� %�� � $hP � $hP ��      >    , ~� �� �� �� �� �� ~� �� ~� ��      >    , �� 	�P "($ 	�P "($ 	� �� 	� �� 	�P      >    , �L :l � :l � F$ �L F$ �L :l      >    , 
�� 	f@ �  	f@ �  	q� 
�� 	q� 
�� 	f@      >    , J0 �8 �( �8 �( � J0 � J0 �8      >    , )��  4� )�  4� )�  @t )��  @t )��  4�      >    , )�P � +�� � +�� �� )�P �� )�P �      >    , ET :l � :l � F$ ET F$ ET :l      >    , 
� :l �( :l �( F$ 
� F$ 
� :l      >    , �� � �( � �( � �� � �� �      >    , g �  �� �  �� ø g ø g �       >    , �� 4 e� 4 e� ?� �� ?� �� 4      >    , � w  �� w  �� �� � �� � w       >    , 	 � �� 
h �� 
h �� 	 � �� 	 � ��      >    , �h !� $d !� $d !�� �h !�� �h !�      >    , &L� � 'g� � 'g� �� &L� �� &L� �      >    , %n �T &�$ �T &�$ � %n � %n �T      >    , #�� � %�� � %�� d #�� d #�� �      >    , �4 H � H � )  �4 )  �4 H      >    , ϐ z� !x\ z� !x\ �X ϐ �X ϐ z�      >    , &�P � )� � )� �X &�P �X &�P �      >    , &�@ 4 'N� 4 'N� ?� &�@ ?� &�@ 4      >    , ~� 0  !b� 0  !b� ;� ~� ;� ~� 0       >    , �4 �@ l �@ l �� �4 �� �4 �@      >    , 	�� !�L 
? !�L 
? !� 	�� !� 	�� !�L      >    , 
7<  � ^   � ^   �� 
7<  �� 
7<  �      >    , �\ Wx 1 Wx 1 c0 �\ c0 �\ Wx      >    , "� �  #�� �  #�� ø "� ø "� �       >    , %�� �� (#d �� (#d �� %�� �� %�� ��      >    , ):� � )� � )� �� ):� �� ):� �      >    , �@ �� T� �� T� �| �@ �| �@ ��      >    , � o� #z o� #z {L � {L � o�      >    , �h �� &� �� &� �� �h �� �h ��      >    , � >4 �L >4 �L I� � I� � >4      >    , �| v� %� v� %� �� �| �� �| v�      >    , &i� !�L 'w� !�L 'w� !� &i� !� &i� !�L      >    , VT ;� <� ;� <� GH VT GH VT ;�      >    , %�p �� )�@ �� )�@ �� %�p �� %�p ��      >    , � � h� � h� �� � �� � �      >    , �0 ', �� ', �� 2� �0 2� �0 ',      >    , (�� |� *<� |� *<� �D (�� �D (�� |�      >    , 
�x O 
�X O 
�X Z� 
�x Z� 
�x O      >    , S� T@ l� T@ l� _� S� _� S� T@      >    , -?� d� .j� d� .j� p� -?� p� -?� d�      >    , )#@ >4 )�8 >4 )�8 I� )#@ I� )#@ >4      >    , +�  �� ,�� �� ,�� �� +�  �� +�  ��      >    , :p �( x� �( x� �� :p �� :p �(      >    , -_<   .;�   .;� � -_< � -_<        >    , $�  d� %T� d� %T� p� $�  p� $�  d�      >    , RL %�L }D %�L }D %� RL %� RL %�L      >    , 
�| �  /$ �  /$ ø 
�| ø 
�| �       >    , d� �4 �� �4 �� �� d� �� d� �4      >    , S� �� � �� � �� S� �� S� ��      >    , �  �� � �� � �D �  �D �  ��      >    , 6` �h e@ �h e@ �  6` �  6` �h      >    , %�h !�L &R� !�L &R� !� %�h !� %�h !�L      >    , "� &l "l� &l "l� &$ "� &$ "� &l      >    , +�� b� -I� b� -I� nX +�� nX +�� b�      >    , (�� �h *�@ �h *�@ �  (�� �  (�� �h      >    , �� �� "�p �� "�p �� �� �� �� ��      >    , "�� Đ "� Đ "� �H "�� �H "�� Đ      >    , �� � �� � �� �� �� �� �� �      >    , �0 eD 
�� eD 
�� p� �0 p� �0 eD      >    , )�� !�L *@ !�L *@ !� )�� !� )�� !�L      >    , \ \ �� \ ��   \   \ \      >    , �� � ^H � ^H � �� � �� �      >    , �p ��   ��   �� �p �� �p ��      >    , �< � �� � �� � �< � �< �      >    , �| 0� E 0� E <d �| <d �| 0�      >    , 9P "b� �� "b� �� "nt 9P "nt 9P "b�      >    , !�< �� $�� �� $�� �� !�< �� !�< ��      >    , �  � ��  � ��  �H �  �H �  �      >    , �� �( ȸ �( ȸ �� �� �� �� �(      >    , �� 	�x -� 	�x -� 	�0 �� 	�0 �� 	�x      >    , � ;� �8 ;� �8 GH � GH � ;�      >    , &�x F� -�$ F� -�$ Rl &�x Rl &�x F�      >    ,  d� ?t  �| ?t  �| K,  d� K,  d� ?t      >    ,  �� 	�x #� 	�x #� 	�0  �� 	�0  �� 	�x      >    , !l� b� !� b� !� nX !l� nX !l� b�      >    , XH  � �  � �  �H XH  �H XH  �      >    , $�| \ %�� \ %��  $�|  $�| \      >    , � =� � =� � I� � I� � =�      >    , �� � � � � �� �� �� �� �      >    , *oH � +܄ � +܄ �� *oH �� *oH �      >    , �� #��  #��  #� �� #� �� #��      >    , �4 $G �� $G �� $R� �4 $R� �4 $G      >    , �� "� �8 "� �8 "�� �� "�� �� "�      >    , �� 	?0 �8 	?0 �8 	J� �� 	J� �� 	?0      >    , �� �$ �� �$ �� �� �� �� �� �$      >    , 3� ~� ߜ ~� ߜ �\ 3� �\ 3� ~�      >    , &� 8T 'b 8T 'b D &� D &� 8T      >    , M�  �X  �  �X  �  � M�  � M�  �X      >    , �x 	� Y� 	� Y� X �x X �x 	�      >    , �� 4 �T 4 �T ?� �� ?� �� 4      >    , G� $�� �x $�� �x $�< G� $�< G� $��      >    , \ � @H � @H �� \ �� \ �      >    , d !=� �� !=� �� !I| d !I| d !=�      >    , #{� >� )<� >� )<� JX #{� JX #{� >�      >    , $�� 	 'b 	 'b 	'� $�� 	'� $�� 	      >    , 
D d� 
�� d� 
�� p� 
D p� 
D d�      >    , � 	� =� 	� =� X � X � 	�      >    , oL ��  4$ ��  4$ � oL � oL ��      >    , �<  !�L  !�L �P �< �P �<       >    , s� �� ' �� ' �| s� �| s� ��      >    , !n� !�< "A� !�< "A� !�� !n� !�� !n� !�<      >    , a� ��  ��  �t a� �t a� ��      >    , �$ �� ct �� ct �t �$ �t �$ ��      >    , 6 !�L �` !�L �` !� 6 !� 6 !�L      >    , �� 	f@ ܌ 	f@ ܌ 	q� �� 	q� �� 	f@      >    , "�� �� #"$ �� #"$ �� "�� �� "�� ��      >    , q� 4P #  4P #  @ q� @ q� 4P      >    , %T #�� & #�� & #�| %T #�| %T #��      >    , �� �, 0� �, 0� �� �� �� �� �,      >    , #� �� 1� �� 1� �L #� �L #� ��      >    , +| �@ ,S� �@ ,S� �� +| �� +| �@      >    , |� ��  �d ��  �d �� |� �� |� ��      >    , '�� (P (�� (P (�� 4 '�� 4 '�� (P      >    , �@ � �  � �  �� �@ �� �@ �      >    , �< i, n� i, n� t� �< t� �< i,      >    , �p S� �� S� �� _� �p _� �p S�      >    , �� �8 eh �8 eh � �� � �� �8      >    , C� eD �  eD �  p� C� p� C� eD      >    , Q 	f@ � 	f@ � 	q� Q 	q� Q 	f@      >    , -�� ld .� ld .� x -�� x -�� ld      >    ,  H �� H �� )   )   H      >    , 
{� >4 � >4 � I� 
{� I� 
{� >4      >    , =� �D �� �D �� �� =� �� =� �D      >    , �� :l 7� :l 7� F$ �� F$ �� :l      >    , )�| F� -�@ F� -�@ Rp )�| Rp )�| F�      >    , ,�p h .@ h .@   ,�p   ,�p h      >    , #�, ";� '3( ";� '3( "Gd #�, "Gd #�, ";�      >    , �� d� T d� T p� �� p� �� d�      >    , �� �  �H �  �H ø �� ø �� �       >    , �d $ � 	V� $ � 	V� $� �d $� �d $ �      >    , 
�� 7� D� 7� D� C< 
�� C< 
�� 7�      >    , < |� (� |� (� �D < �D < |�      >    , � |� 0 |� 0 �D � �D � |�      >    , �   �(   �(  � �  � �       >    , ,�� :l -(� :l -(� F$ ,�� F$ ,�� :l      >    , j� �� r �� r �� j� �� j� ��      >    , :$ 
ɸ  ]( 
ɸ  ]( 
�p :$ 
�p :$ 
ɸ      >    , � >4 �( >4 �( I� � I� � >4      >    ,  f�  �X #��  �X #��  �  f�  �  f�  �X      >    ,  @  � ��  � ��  �H  @  �H  @  �      >    , (8� !�\ )B� !�\ )B� " (8� " (8� !�\      >    , %�X � &�� � &�� �� %�X �� %�X �      >    , � �� �� �� �� �� � �� � ��      >    , � $ L $ L "� � "� � $      >    , #�  �8 $L� �8 $L� � #�  � #�  �8      >    , )�0 4 *�8 4 *�8 ?� )�0 ?� )�0 4      >    , H< ٜ �� ٜ �� �T H< �T H< ٜ      >    , Լ �� O� �� O� �H Լ �H Լ ��      >    , U� �� b� �� b� | U� | U� ��      >    , @ H M  H M  )  @ )  @ H      >    , Ah 	�� p  	�� p  
h Ah 
h Ah 	��      >    , � :l � :l � F$ � F$ � :l      >    , *4� H *ܨ H *ܨ )  *4� )  *4� H      >    , �(   >�   >� � �( � �(        >    , +4 i� , i� , u� +4 u� +4 i�      >    , MH #�� pL #�� pL #� MH #� MH #��      >    , hT �( �� �( �� �� hT �� hT �(      >    , %R� d� %�� d� %�� p� %R� p� %R� d�      >    , � �� �� �� �� �� � �� � ��      >    , �� C a\ C a\ N� �� N� �� C      >    , .P �� -� �� -� �� .P �� .P ��      >    , & � F� (N\ F� (N\ Rp & � Rp & � F�      >    ,  x� �h  �< �h  �< �   x� �   x� �h      >    , -� �� -M� �� -M� �t -� �t -� ��      >    , !� �8 X� �8 X� �� !� �� !� �8      >    , � 	�P �h 	�P �h 	� � 	� � 	�P      >    , z� �| �� �| �� �4 z� �4 z� �|      >    , $հ �( %`\ �( %`\ �� $հ �� $հ �(      >    , { 
�P 2� 
�P 2� 
� { 
� { 
�P      >    , *>t �� ,6\ �� ,6\ �� *>t �� *>t ��      >    , +�� �D ,�� �D ,�� �� +�� �� +�� �D      >    , m� � w@ � w@ �� m� �� m� �      >    , ~<  �� �  �� �  �8 ~<  �8 ~<  ��      >    , -�  �� �h  �� �h  �8 -�  �8 -�  ��      >    , %�D #�� &� #�� &� #� %�D #� %�D #��      >    , (g� d� *� d� *� pl (g� pl (g� d�      >    , )�l 	�� *4 	�� *4 
� )�l 
� )�l 	��      >    , 	�� � 
�( � 
�( �� 	�� �� 	�� �      >    , 	�� � Z@ � Z@ �� 	�� �� 	�� �      >    , (, !G� W !G� W !S@ (, !S@ (, !G�      >    , ר �( j$ �( j$ �� ר �� ר �(      >    , 3� b� �( b� �( nX 3� nX 3� b�      >    , $�X '@� $�8 '@� $�8 'L� $�X 'L� $�X '@�      >    , %%� %�  %P� %�  %P� %�� %%� %�� %%� %�       >    , u( �� :l �� :l �T u( �T u( ��      >    , �< O� F� O� F� [� �< [� �< O�      >    , q  �  �� �  �� ø q  ø q  �       >    , i0 � ( � ( � i0 � i0 �      >    , }� $ �� $ �� "� }� "� }� $      >    , X� � �� � �� �� X� �� X� �      >    ,  0< Đ  �� Đ  �� �H  0< �H  0< Đ      >    , !�� �� "l �� "l �� !�� �� !�� ��      >    , ct hT �d hT �d t ct t ct hT      >    , �L #�� �8 #�� �8 $� �L $� �L #��      >    , �4 %�L � %�L � %� �4 %� �4 %�L      >    , 
�P &J� �, &J� �, &Vt 
�P &Vt 
�P &J�      >    , Ҩ d� I� d� I� p� Ҩ p� Ҩ d�      >    , ?T #�� 	� #�� 	� #� ?T #� ?T #��      >    , ?T !� �8 !� �8 !�� ?T !�� ?T !�      >    , `� �� �T �� �T �T `� �T `� ��      >    , (�� � )�� � )��  � (��  � (�� �      >    , (� %�d +d %�d +d %� (� %� (� %�d      >    , � �� � �� � �D � �D � ��      >    , �� %�\ �� %�\ �� %� �� %� �� %�\      >    , �| � �� � �� �� �| �� �| �      >    , �h �T '0 �T '0 � �h � �h �T      >    , � �X � �X � � � � � �X      >    , �< �$ �x �$ �x �� �< �� �< �$      >    , :� "� �� "� �� "�� :� "�� :� "�      >    , �D �� & �� & �| �D �| �D ��      >    , �( �� Gl �� Gl �| �( �| �( ��      >    , �p !�< � !�< � !�� �p !�� �p !�<      >    , B� $ �� $ �� "� B� "� B� $      >    , 	�� #�� 
�� #�� 
�� #� 	�� #� 	�� #��      >    , M  ;� L� ;� L� GH M  GH M  ;�      >    , Sh �� � �� � �� Sh �� Sh ��      >    , �L %�\ ( %�\ ( %� �L %� �L %�\      >    , 	N� #�� m� #�� m� $� 	N� $� 	N� #��      >    , ʌ �D � �D � �� ʌ �� ʌ �D      >    , &  �� )V �� )V � &  � &  ��      >    , 4 �� _d �� _d �� 4 �� 4 ��      >    , �h 4 �0 4 �0 ?� �h ?� �h 4      >    , 'e� ', )e� ', )e� 2� 'e� 2� 'e� ',      >    , �0 b� _  b� _  nX �0 nX �0 b�      >    , �� ʬ *� ʬ *� �d �� �d �� ʬ      >    , 	�� "�� �� "�� �� "�� 	�� "�� 	�� "��      >    , *� �8 *�� �8 *�� � *� � *� �8      >    , *@ 	 +q 	 +q � *@ � *@ 	      >    , 	�h �� 
3T �� 
3T �D 	�h �D 	�h ��      >    , &�$ �� '#� �� '#� 	� &�$ 	� &�$ ��      >    , �@ JT Ҁ JT Ҁ V �@ V �@ JT      >    , v� �� >� �� >� �t v� �t v� ��      >    , #CX �D $dh �D $dh �� #CX �� #CX �D      >    , a� 7� �� 7� �� C< a� C< a� 7�      >    , @( !�L �L !�L �L !� @( !� @( !�L      >    , ,� �� ,� �� ,� �D ,� �D ,� ��      >    , �< � h � h �� �< �� �< �      >    , -0 	f@ !T 	f@ !T 	q� -0 	q� -0 	f@      >    , �H �� �� �� �� �| �H �| �H ��      >    , .p �L � �L � � .p � .p �L      >    , '�  i� ($ i� ($ u� '�  u� '�  i�      >    , %T �( %�� �( %�� �� %T �� %T �(      >    , q@ �( 8x �( 8x �� q@ �� q@ �(      >    , �� x� C� x� C� �\ �� �\ �� x�      >    , \� #�� �� #�� �� #� \� #� \� #��      >    , 	q� i� 
s� i� 
s� u� 	q� u� 	q� i�      >    ,  A� H !� H !� )   A� )   A� H      >    , <� ;� ip ;� ip GH <� GH <� ;�      >    , %< >4 V >4 V I� %< I� %< >4      >    , '�l � )�� � )��  8 '�l  8 '�l �      >    , .� ;� .j� ;� .j� GH .� GH .� ;�      >    , )� d� �� d� �� pl )� pl )� d�      >    , '0 � �� � �� @ '0 @ '0 �      >    , �� � 	� � 	� � �� � �� �      >    , 8 4 l 4 l ?� 8 ?� 8 4      >    , �< �D a� �D a� �� �< �� �< �D      >    , � ٜ Ex ٜ Ex �T � �T � ٜ      >    , |� �D ?� �D ?� �� |� �� |� �D      >    , wD 4 �8 4 �8 %� wD %� wD 4      >    , �  �� S$  �� S$  �8 �  �8 �  ��      >    , � Z� �  Z� �  fd � fd � Z�      >    , (+4 �� *% �� *% �� (+4 �� (+4 ��      >    , +� d� -( d� -( pl +� pl +� d�      >    , "� �� �@ �� �@ �� "� �� "� ��      >    , �X �� h �� h �t �X �t �X ��      >    , ��   �x   �x � �� � ��        >    , �h ��  v� ��  v� �| �h �| �h ��      >    , �D #�� i, #�� i, #�| �D #�| �D #��      >    , �| �� � �� � �� �| �� �| ��      >    , *�� 	f@ +�� 	f@ +�� 	q� *�� 	q� *�� 	f@      >    , -�� �� .S` �� .S` �� -�� �� -�� ��      >    , }� b� !�$ b� !�$ nT }� nT }� b�      >    , Ѩ 	�8 s� 	�8 s� 	�� Ѩ 	�� Ѩ 	�8      >    , ,� O �� O �� Z� ,� Z� ,� O      >    , x< ?t �� ?t �� K, x< K, x< ?t      >    , �� t � t � , �� , �� t      >    , E� Z� x` Z� x` fd E� fd E� Z�      >    , �� � X� � X�  8 ��  8 �� �      >    ,  � #�� !G� #�� !G� #�|  � #�|  � #��      >    , � !�L �� !�L �� !� � !� � !�L      >    , �� i� �@ i� �@ u� �� u� �� i�      >    , ;  ~@ j  ~@ j  �� ;  �� ;  ~@      >    , #�\  � $�   � $�   �H #�\  �H #�\  �      >    , tx �X � �X � � tx � tx �X      >    , f� eD f� eD f� p� f� p� f� eD      >    , P0 �T �� �T �� � P0 � P0 �T      >    , '�� !�< )| !�< )| !�� '�� !�� '�� !�<      >    , �� ~@ <@ ~@ <@ �� �� �� �� ~@      >    , �\ � h � h � �\ � �\ �      >    , :� d� <� d� <� pL :� pL :� d�      >    , *[� �( +"� �( +"� �� *[� �� *[� �(      >    , �� � �� � �� � �� � �� �      >    , - � �P -t� �P -t� � - � � - � �P      >    , !C� �P !r� �P !r� � !C� � !C� �P      >    , k� �� �� �� �� l k� l k� ��      >    , �� |� r� |� r� �D �� �D �� |�      >    , -Є 	j( -�d 	j( -�d 	u� -Є 	u� -Є 	j(      >    , ^l %�\ @ %�\ @ %� ^l %� ^l %�\      >    , ~� !(H �$ !(H �$ !4  ~� !4  ~� !(H      >    , 	Ѭ \ m� \ m�   	Ѭ   	Ѭ \      >    , +<\ \ ,cH \ ,cH  +<\  +<\ \      >    , ,aT \ -�h \ -�h  ,aT  ,aT \      >    , S� �\ @ �\ @ � S� � S� �\      >    , #f� &1X )�� &1X )�� &= #f� &= #f� &1X      >    , ( =�  =�  I� ( I� ( =�      >    , x �� � �� � �� x �� x ��      >    , �l � 5h � 5h � �l � �l �      >    , 'Pt `< '�� `< '�� k� 'Pt k� 'Pt `<      >    , 9� |� Z� |� Z� �D 9� �D 9� |�      >    , � �T � �T � � � � � �T      >    , �� ʬ !Ĉ ʬ !Ĉ �d �� �d �� ʬ      >    , �� �l h� �l h� �$ �� �$ �� �l      >    , X� eD �P eD �P p� X� p� X� eD      >    , �� 4� ۔ 4� ۔ @L �� @L �� 4�      >    , !� 0� $�� 0� $�� <d !� <d !� 0�      >    , 	�L %�\ 
k� %�\ 
k� %� 	�L %� 	�L %�\      >    , l� %�L �$ %�L �$ %� l� %� l� %�L      >    , �   �(   �( � � � �        >    , ¼ Wx  d Wx  d c0 ¼ c0 ¼ Wx      >    , 5  	� X$ 	� X$ X 5  X 5  	�      >    , �� 4P �� 4P �� @ �� @ �� 4P      >    , 	�� 
� �D 
� �D 
%� 	�� 
%� 	�� 
�      >    , &� �0 �� �0 �� �� &� �� &� �0      >    , 	'� � 
)� � 
)� �� 	'� �� 	'� �      >    , �\ [ Ƥ [ Ƥ f� �\ f� �\ [      >    , � !`� �� !`� �� !l� � !l� � !`�      >    , "�� �� "� �� "� �� "�� �� "�� ��      >    , μ L a8 L a8 ( μ ( μ L      >    , {� � 	�d � 	�d �� {� �� {� �      >    , )  �� )�� �� )�� �| )  �| )  ��      >    , �\  � ��  � ��  �H �\  �H �\  �      >    , 
�t �� �` �� �` �� 
�t �� 
�t ��      >    , � �$ 
, �$ 
, � � � � �$      >    , `� �� �� �� �� �T `� �T `� ��      >    , h� =� �h =� �h I� h� I� h� =�      >    , �� � Sl � Sl �� �� �� �� �      >    , qh � 6� � 6� �� qh �� qh �      >    , VX e� x e� x qh VX qh VX e�      >    , � >� �� >� �� JX � JX � >�      >    , N� F� F$ F� F$ Rp N� Rp N� F�      >    , �l [ h [ h f� �l f� �l [      >    , � d� 7� d� 7� p� � p� � d�      >    , 	�� 	�P �� 	�P �� 	� 	�� 	� 	�� 	�P      >    , �T �� �� �� �� �� �T �� �T ��      >    ,  �� �� �� �� �|  �|  ��      >    , $�| ٜ &9( ٜ &9( �T $�| �T $�| ٜ      >    , � �$ � �$ � � � � � �$      >    , !�� d� "j� d� "j� p� !�� p� !�� d�      >    , +H 4 ,� 4 ,� ?� +H ?� +H 4      >    , M� �|  �� �|  �� �4 M� �4 M� �|      >    , +� �4 +4� �4 +4� �� +� �� +� �4      >    , ,�  #�� -x� #�� -x� #� ,�  #� ,�  #��      >    , +q 7� +�� 7� +�� C\ +q C\ +q 7�      >    , �� �(  � �(  � �� �� �� �� �(      >    , -p� #�� .� #�� .� $� -p� $� -p� #��      >    , �d &�� m� &�� m� 'T �d 'T �d &��      >    , }� 4 	G  4 	G  ?� }� ?� }� 4      >    , 
T� �� m� �� m� �| 
T� �| 
T� ��      >    , (� >4 eh >4 eh I� (� I� (� >4      >    , � 	�P J 	�P J 	� � 	� � 	�P      >    , � �� Px �� Px �@ � �@ � ��      >    , �0 ٜ � ٜ � �T �0 �T �0 ٜ      >    , !� !�L #(  !�L #(  !� !� !� !� !�L      >    , T� �� �D �� �D �D T� �D T� ��      >    , �� �� | �� | �D �� �D �� ��      >    , $� 4 %׀ 4 %׀ ?� $� ?� $� 4      >    , �� 4 �� 4 �� ?� �� ?� �� 4      >    , (�� �  )�H �  )�H ø (�� ø (�� �       >    , '�\ ;� (�  ;� (�  GH '�\ GH '�\ ;�      >    , | �, � �, � �� | �� | �,      >    , �h 4P E 4P E @ �h @ �h 4P      >    , �<   9P   9P � �< � �<        >    , 	�h 
�� 
�D 
�� 
�D \ 	�h \ 	�h 
��      >    , !�� :l "�  :l "�  F$ !�� F$ !�� :l      >    , �4 �T �� �T �� � �4 � �4 �T      >    , W� ֌ �x ֌ �x �D W� �D W� ֌      >    , hT �l �4 �l �4 �$ hT �$ hT �l      >    , �� z� =� z� =� �� �� �� �� z�      >    , 	�H ٜ 	�( ٜ 	�( �T 	�H �T 	�H ٜ      >    , �( �\ 2� �\ 2� � �( � �( �\      >    , ' �T � �T � � ' � ' �T      >    , *_� �` *� �` *� � *_� � *_� �`      >    , � L ^ L ^  �  � L      >    , Q, 
`@ @ 
`@ @ 
k� Q, 
k� Q, 
`@      >    , .X �  .08 �  .08 ø .X ø .X �       >    , )a� � *(� � *(� �� )a� �� )a� �      >    , �� �( "x8 �( "x8 �� �� �� �� �(      >    , .� �D O� �D O� �� .� �� .� �D      >    , Z� � [� � [� �� Z� �� Z� �      >    , k� �� RL �� RL �| k� �| k� ��      >    , .&t �� .UT �� .UT �� .&t �� .&t ��      >    , �0 f< �l f< �l q� �0 q� �0 f<      >    , s� �� �` �� �` � s� � s� ��      >    , WT �� �4 �� �4 ڔ WT ڔ WT ��      >    , #� �( $p  �( $p  �� #� �� #� �(      >    , �\ 
= y� 
= y� 
H� �\ 
H� �\ 
=      >    , 
^L 	bX 
�, 	bX 
�, 	n 
^L 	n 
^L 	bX      >    , �� &'� GH &'� GH &3L �� &3L �� &'�      >    , (� � )�  � )�  �� (� �� (� �      >    , �$  �� ;�  �� ;�  �8 �$  �8 �$  ��      >    , , i� ,�  i� ,�  u� , u� , i�      >    , s4 	�P �H 	�P �H 	� s4 	� s4 	�P      >    , � !�L 18 !�L 18 !� � !� � !�L      >    , .� �� 0� �� 0� �D .� �D .� ��      >    , (�� �� ) �� ) �| (�� �| (�� ��      >    , 2X 4P �x 4P �x @ 2X @ 2X 4P      >    , � ;� �� ;� �� GH � GH � ;�      >    , � H � H � )  � )  � H      >    , ֈ �d h �d h � ֈ � ֈ �d      >    , Z �| {( �| {( �4 Z �4 Z �|      >    , � �, l` �, l` �� � �� � �,      >    , G$ �� n� �� n� �� G$ �� G$ ��      >    , 4 4P �� 4P �� @ 4 @ 4 4P      >    , � �� �� �� �� �� � �� � ��      >    , �  �� "� �� "� �L �  �L �  ��      >    ,  A� ^l 1� ^l 1� j$  A� j$  A� ^l      >    , (� 	f@ )�` 	f@ )�` 	q� (� 	q� (� 	f@      >    , a| #�� p� #�� p� #�| a| #�| a| #��      >    , !� � "M@ � "M@ �� !� �� !� �      >    , < ;� r� ;� r� GH < GH < ;�      >    , �h zX  zX  � �h � �h zX      >    ,   �� �(  �� �(  �x   �x   ��      >    , "�� �8 #�� �8 #�� � "�� � "�� �8      >    , v� �4 �\ �4 �\ �� v� �� v� �4      >    , B@ :l �� :l �� F$ B@ F$ B@ :l      >    , ,Ԑ d� -(� d� -(� p� ,Ԑ p� ,Ԑ d�      >    , �� m| e@ m| e@ y4 �� y4 �� m|      >    , M� �� |� �� |� �D M� �D M� ��      >    , 9 d� %` d� %` p� 9 p� 9 d�      >    , c �8 �� �8 �� � c � c �8      >    , -�@ �� .08 �� .08 �| -�@ �| -�@ ��      >    ,   hT ~� hT ~� t   t   hT      >    , (e� d� ) d� ) p� (e� p� (e� d�      >    , �� �� 	x �� 	x �� �� �� �� ��      >    , �� 	f@ �T 	f@ �T 	q� �� 	q� �� 	f@      >    , #CX %�  #r8 %�  #r8 %�� #CX %�� #CX %�       >    ,  �t :l !&T :l !&T F$  �t F$  �t :l      >    ,  �t JT %$ JT %$ V  �t V  �t JT      >    , �� H � H � )  �� )  �� H      >    , .( 4 Č 4 Č ?� .( ?� .( 4      >    , h "� R  "� R  "$< h "$< h "�      >    , 'i� �� '�P �� '�P �� 'i� �� 'i� ��      >    , )>� SH +� SH +� _  )>� _  )>� SH      >    , 
� � 
L� � 
L� %� 
� %� 
� �      >    , "� 	?0 #5� 	?0 #5� 	J� "� 	J� "� 	?0      >    , #5� � $
� � $
� �� #5� �� #5� �      >    , �P g� -�@ g� -�@ s� �P s� �P g�      >    , �� !�\ �� !�\ �� " �� " �� !�\      >    , �t H �� H �� )  �t )  �t H      >    , �P l< �p l< �p w� �P w� �P l<      >    , i0 |� �p |� �p �D i0 �D i0 |�      >    , �� >T �� >T �� J �� J �� >T      >    , �� 	�P �h 	�P �h 	� �� 	� �� 	�P      >    , S� ET �d ET �d Q S� Q S� ET      >    , �| 	?0 !W( 	?0 !W( 	J� �| 	J� �| 	?0      >    , qh $ � $ � "� qh "� qh $      >    , �t �8 u, �8 u, � �t � �t �8      >    , � �8 � �8 � � � � � �8      >    , � �( �� �( �� �� � �� � �(      >    , �4 !�< 	�d !�< 	�d !�� �4 !�� �4 !�<      >    , "5� \ #M \ #M  "5�  "5� \      >    , � |� ;� |� ;� �D � �D � |�      >    , � � � � � (L � (L � �      >    , p� z� �� z� �� �X p� �X p� z�      >    ,  �� �� !� �� !� ��  �� ��  �� ��      >    , � 4 �h 4 �h ?� � ?� � 4      >    ,    	�x  =� 	�x  =� 	�0    	�0    	�x      >    , %y� � &@� � &@� �� %y� �� %y� �      >    , �T %�L #� %�L #� %� �T %� �T %�L      >    , �� �D 
8 �D 
8 �� �� �� �� �D      >    , � 4 �( 4 �( ?� � ?� � 4      >    , ϐ #�� � #�� � #�| ϐ #�| ϐ #��      >    , }� #�� �� #�� �� #� }� #� }� #��      >    , ,�8 �� -p� �� -p� �| ,�8 �| ,�8 ��      >    , #� ȼ #�� ȼ #�� �t #� �t #� ȼ      >    , �| �  {( �  {( ø �| ø �| �       >    , 8 !�L �L !�L �L !� 8 !� 8 !�L      >    , 
�| t 8 t 8 , 
�| , 
�| t      >    , �@ $f\ �  $f\ �  $r �@ $r �@ $f\      >    , � �� ˨ �� ˨ �H � �H � ��      >    , � b� 	;H b� 	;H nX � nX � b�      >    , -�� #�� .E� #�� .E� #� -�� #� -�� #��      >    ,  #�� :� #�� :� #�  #�  #��      >    , ,G� � .� � .� �� ,G� �� ,G� �      >    , k� �� �\ �� �\ �@ k� �@ k� ��      >    , "d� 	 $�� 	 $�� 	'� "d� 	'� "d� 	      >    , � 0� 	�� 0� 	�� <d � <d � 0�      >    , � :l ! :l ! F$ � F$ � :l      >    , �� %�L �\ %�L �\ %� �� %� �� %�L      >    , *,� �D +x� �D +x� �� *,� �� *,� �D      >    , $�D � %� � %� �� $�D �� $�D �      >    , "�� = '0 = '0 H� "�� H� "�� =      >    , .S` �� .�4 �� .�4 ֬ .S` ֬ .S` ��      >    , 1 >4 \ >4 \ I� 1 I� 1 >4      >    , 
� b� -� b� -� nT 
� nT 
� b�      >    , .( �� �l �� �l �D .( �D .( ��      >    , #�� �� $%� �� $%� �L #�� �L #�� ��      >    , � [| @ [| @ g4 � g4 � [|      >    , Z� ^� 
�� ^� 
�� jL Z� jL Z� ^�      >    , D � ^� � ^� +� D +� D �      >    , �� :l |� :l |� F$ �� F$ �� :l      >    , $�h �� %C �� %C �� $�h �� $�h ��      >    , &| �| �� �| �� �4 &| �4 &| �|      >    , �l >4 �` >4 �` I� �l I� �l >4      >    , �� � �� � �� �� �� �� �� �      >    , 	� �D 8� �D 8� �� 	� �� 	� �D      >    , 
h L 
�x L 
�x ( 
h ( 
h L      >    , H@ 
= ܌ 
= ܌ 
H� H@ 
H� H@ 
=      >    , �  � |L  � |L d � d �  �      >    , � $ !	 $ !	 "� � "� � $      >    , "5� �| #�d �| #�d �4 "5� �4 "5� �|      >    ,  _ � !� � !�  8  _  8  _ �      >    ,  � �P !"l �P !"l �  � �  � �P      >    ,  �4 
�l �4 
�l ��  ��  �4      >    , #K( ?t &o� ?t &o� K, #K( K, #K( ?t      >    , ,� ', .�( ', .�( 2� ,� 2� ,� ',      >    , 	� �8 ؠ �8 ؠ � 	� � 	� �8      >    , )h �T �  �T �  � )h � )h �T      >    , �� = 	� = 	� H� �� H� �� =      >    , �� �8 �L �8 �L � �� � �� �8      >    , 
  � 
T� � 
T� �� 
  �� 
  �      >    , �  u0 �$  u0 �$  �� �  �� �  u0      >    , �� >4 �` >4 �` I� �� I� �� >4      >    , !, _� '/@ _� '/@ kH !, kH !, _�      >    , �` b� �@ b� �@ n� �` n� �` b�      >    , I� &'� V� &'� V� &3L I� &3L I� &'�      >    , �, #�� �8 #�� �8 #� �, #� �, #��      >    , �L �� �� �� �� �T �L �T �L ��      >    ,   �� (p �� (p �T   �T   ��      >    , � 7�  *` 7�  *` C< � C< � 7�      >    , &  ȼ '�� ȼ '�� �t &  �t &  ȼ      >    , R� �� 5h �� 5h �| R� �| R� ��      >    , 	�p H �@ H �@ )  	�p )  	�p H      >    , (]� G� )Fh G� )Fh SH (]� SH (]� G�      >    , �| !�\ �� !�\ �� " �| " �| !�\      >    , �T %�\ �� %�\ �� %� �T %� �T %�\      >    , 0� v� cP v� cP �� 0� �� 0� v�      >    , � ,� &4 ,� &4 8� � 8� � ,�      >    , &� :l 'ð :l 'ð F$ &� F$ &� :l      >    , �\ A� �� A� �� MD �\ MD �\ A�      >    , 	�P &l 
D� &l 
D� &$ 	�P &$ 	�P &l      >    , �L �\ 	;H �\ 	;H � �L � �L �\      >    , 4  �� �  �� �  �8 4  �8 4  ��      >    , #� "^� %^h "^� %^h "j� #� "j� #� "^�      >    , 
( 	f@ -, 	f@ -, 	q� 
( 	q� 
( 	f@      >    , '�X $� (�� $� (�� $x '�X $x '�X $�      >    , )LD #�� +d #�� +d #� )LD #� )LD #��      >    , (P ٜ Y$ ٜ Y$ �T (P �T (P ٜ      >    , �L !� �� !� �� !�� �L !�� �L !�      >    , )�T 	� *B\ 	� *B\ X )�T X )�T 	�      >    , $հ %�  %-� %�  %-� %�� $հ %�� $հ %�       >    , l� �� ȸ �� ȸ �l l� �l l� ��      >    , 	D �� 
� �� 
� �T 	D �T 	D ��      >    , {L �T � �T � � {L � {L �T      >    , '�  
� '�� 
� '�� � '�  � '�  
�      >    ,  � � !S@ � !S@ ��  � ��  � �      >    , )�X  � )��  � )��  d )�X  d )�X  �      >    , )� _� *� _� *� kH )� kH )� _�      >    , !C� �� !�( �� !�( �� !C� �� !C� ��      >    , ,�� #� -�h #� -�h /H ,�� /H ,�� #�      >    , +m0 �( ,�d �( ,�d �� +m0 �� +m0 �(      >    , �� "�� �� "�� �� "�� �� "�� �� "��      >    , g �T �T �T �T � g � g �T      >    , '�  � (F� � (F� �� '�  �� '�  �      >    , (D� � )#@ � )#@ �� (D� �� (D� �      >    , �P �< � �< � �� �P �� �P �<      >    , �\ 4 |  4 |  ?� �\ ?� �\ 4      >    , "�� d� $`� d� $`� p� "�� p� "�� d�      >    , ߠ 6� �� 6� �� B� ߠ B� ߠ 6�      >    , �� � Đ � Đ � �� � �� �      >    , H m| Y� m| Y� y4 H y4 H m|      >    , "�\ !�\ ${� !�\ ${� " "�\ " "�\ !�\      >    , �h �� x� �� x� �T �h �T �h ��      >    , �X �� �\ �� �\ �T �X �T �X ��      >    , � , ;h , ;h  � �  � � ,      >    , � �8 � �8 � � � � � �8      >    , ��  d ��  d ��  ��  ��  d      >    , w !�< F$ !�< F$ !�� w !�� w !�<      >    , % !�L %�� !�L %�� !� % !� % !�L      >    , -�� ET -�d ET -�d Q -�� Q -�� ET      >    , $�  �� $�� �� $�� �l $�  �l $�  ��      >    , %�� ~@ &3L ~@ &3L �� %�� �� %�� ~@      >    , 
�| �� b �� b �T 
�| �T 
�| ��      >    , $L� 
� $w� 
� $w� � $L� � $L� 
�      >    , �� $ +� $ +� "� �� "� �� $      >    , (X  <h *�� <h *�� H  (X  H  (X  <h      >    , AD 
�x �d 
�x �d 
�0 AD 
�0 AD 
�x      >    , �  � �  � �  � �  � �  �      >    , |� hT  hT  t |� t |� hT      >    , &�� d� '�� d� '�� pl &�� pl &�� d�      >    , �� �� h �� h �D �� �D �� ��      >    , :� �l qD �l qD $ :� $ :� �l      >    , �P �4 \ �4 \ �� �P �� �P �4      >    , X$ �� ,�x �� ,�x ڔ X$ ڔ X$ ��      >    , $X� d� $�� d� $�� p� $X� p� $X� d�      >    , �8 �� � �� � �� �8 �� �8 ��      >    , �< � �� � �� �� �< �� �< �      >    ,  � � !�\ � !�\ ��  � ��  � �      >    , $�� �� &� �� &� �| $�� �| $�� ��      >    , L( �� M� �� M� �T L( �T L( ��      >    , +�X !�< ,�h !�< ,�h !�� +�X !�� +�X !�<      >    , :p #�� �@ #�� �@ $� :p $� :p #��      >    , �H ]� ( ]� ( iL �H iL �H ]�      >    , 	�� � �h � �h �L 	�� �L 	�� �      >    , �L 
�h 5h 
�h 5h 
�  �L 
�  �L 
�h      >    , &�P � (�p � (�p �8 &�P �8 &�P �      >    , Ԙ 	�P �� 	�P �� 	� Ԙ 	� Ԙ 	�P      >    , !=� !�L !� !�L !� !� !=� !� !=� !�L      >    , *ڴ !�\ +@ !�\ +@ " *ڴ " *ڴ !�\      >    ,    ��  :  ��  :  ��    ��    ��      >    , 
� �� �� �� �� �D 
� �D 
� ��      >    , � a� �� a� �� m� � m� � a�      >    , �� �� �� �� �� �� �� �� �� ��      >    , X� 
`@ � 
`@ � 
k� X� 
k� X� 
`@      >    , P a| q  a| q  m4 P m4 P a|      >    , " T m| $�� m| $�� y4 " T y4 " T m|      >    , @ ,� �� ,� �� 8� @ 8� @ ,�      >    , �� ,� P� ,� P� 8� �� 8� �� ,�      >    , 0�  �� 0�  �� 0�  �8 0�  �8 0�  ��      >    , !� �� )<� �� )<� �� !� �� !� ��      >    , ,k �4 ,�� �4 ,�� �� ,k �� ,k �4      >    , $� >4 �� >4 �� I� $� I� $� >4      >    , �  v� !�� v� !�� �� �  �� �  v�      >    , � �  Bd �  Bd ø � ø � �       >    , �� \ �� \ ��  ��  �� \      >    , 6 #�� �� #�� �� #� 6 #� 6 #��      >    , '< 	bX '�� 	bX '�� 	n '< 	n '< 	bX      >    , %=4 X &� X &� ! %=4 ! %=4 X      >    , �| !�L �0 !�L �0 !� �| !� �| !�L      >    , �D Yd �d Yd �d e �D e �D Yd      >    , �� s �� s �� ~� �� ~� �� s      >    , !�� �� #d� �� #d� �D !�� �D !�� ��      >    ,  6 � %׀ � %׀ ��  6 ��  6 �      >    , $9p �\ 'H �\ 'H � $9p � $9p �\      >    , '�P � (�� � (�� �� '�P �� '�P �      >    , )�� &l ,� &l ,� &$ )�� &$ )�� &l      >    , % 	f@ ' 	f@ ' 	q� % 	q� % 	f@      >    , +8 	f@ <� 	f@ <� 	q� +8 	q� +8 	f@      >    , #^� � $$ � $$ �� #^� �� #^� �      >    , 
V| 0� 	� 0� 	� <h 
V| <h 
V| 0�      >    , �( �  ?� �  ?� � �( � �( �      >    , � �T 7� �T 7� � � � � �T      >    , ,( ;� ,�� ;� ,�� GH ,( GH ,( ;�      >    , ֐ � �� � �� �� ֐ �� ֐ �      >    ,  6 %�\ !� %�\ !� %�  6 %�  6 %�\      >    , )�X {� *J, {� *J, �� )�X �� )�X {�      >    , �� %$ l< %$ l< %!� �� %!� �� %$      >    , �@ Z� �( Z� �( fd �@ fd �@ Z�      >    , (� �� *B\ �� *B\ �� (� �� (� ��      >    , 'T �� �h �� �h �� 'T �� 'T ��      >    , � "l d "l d "($ � "($ � "l      >    ,  O| >4 !,0 >4 !,0 I�  O| I�  O| >4      >    , !&T $ #� $ #� "� !&T "� !&T $      >    , � �� 28 �� 28 �T � �T � ��      >    , `� :l � :l � F$ `� F$ `� :l      >    , � � �d � �d �� � �� � �      >    , c� � �( � �( �� c� �� c� �      >    , �t b� �L b� �L nX �t nX �t b�      >    , �D @l �$ @l �$ L$ �D L$ �D @l      >    , '� �� )	� �� )	� �� '� �� '� ��      >    , O� �T Ҥ �T Ҥ � O� � O� �T      >    , )�� #�� -E� #�� -E� $� )�� $� )�� #��      >    , +� ~� �X ~� �X �\ +� �\ +� ~�      >    , (/  �� )V  �� )V  �8 (/  �8 (/  ��      >    ,   �P %y� �P %y�       �P      >    , � �� ` �� ` �D � �D � ��      >    , � a� [8 a� [8 m� � m� � a�      >    , �� !�< � !�< � !�� �� !�� �� !�<      >    , 	�0 f< 8 f< 8 q� 	�0 q� 	�0 f<      >    , X  � �@  � �@  �H X  �H X  �      >    , !b�  �� "j�  �� "j�  �8 !b�  �8 !b�  ��      >    , 
 !�L 8� !�L 8� !� 
 !� 
 !�L      >    , 8x �� I� �� I� �| 8x �| 8x ��      >    , �� �� �x �� �x �t �� �t �� ��      >    , .L x ], x ], '0 .L '0 .L x      >    , )�� �� -@ �� -@ �� )�� �� )�� ��      >    , 4� � �� � �� �� 4� �� 4� �      >    , }h G� 
 G� 
 S� }h S� }h G�      >    , !j� x� ".  x� ".  �\ !j� �\ !j� x�      >    , �| ̤ ڸ ̤ ڸ �\ �| �\ �| ̤      >    , "j� �T "� �T "� � "j� � "j� �T      >    , 
p $�� �l $�� �l $�� 
p $�� 
p $��      >    , +K� �4 +�� �4 +�� �� +K� �� +K� �4      >    , +� i� )� i� )� u� +� u� +� i�      >    , �| �� �x �� �x �� �| �� �| ��      >    , ;l �L 	l �L 	l � ;l � ;l �L      >    , �\ L +]� L +]� ( �\ ( �\ L      >    , !  =� "� =� "� I� !  I� !  =�      >    , �0 �� e �� e �t �0 �t �0 ��      >    , �� 	�P P 	�P P 	� �� 	� �� 	�P      >    ,  | �  d� �  d� ø  | ø  | �       >    , H< �� �$ �� �$ �| H< �| H< ��      >    , � S� \� S� \� _� � _� � S�      >    , �| �� 
'� �� 
'� �� �| �� �| ��      >    , (� i� ){$ i� ){$ u� (� u� (� i�      >    , �h 	� <� 	� <� X �h X �h 	�      >    , "� � #z � #z �� "� �� "� �      >    , �� 4  � 4  � ?� �� ?� �� 4      >    , � �P @ �P @ � � � � �P      >    , �h �� @ �� @ �� �h �� �h ��      >    , /� �t �d �t �d �, /� �, /� �t      >    , $�X &0 '�@ &0 '�@ &� $�X &� $�X &0      >    , &р  � '�<  � '�< � &р � &р  �      >    , � &l RH &l RH &$ � &$ � &l      >    , ڼ � cP � cP �p ڼ �p ڼ �      >    , %� o, '3( o, '3( z� %� z� %� o,      >    , ְ >4 �` >4 �` I� ְ I� ְ >4      >    , I� � �d � �d �� I� �� I� �      >    , $� 	�� `� 	�� `� 
� $� 
� $� 	��      >    , �| 
� | 
� | 
%� �| 
%� �| 
�      >    , '�L �� (Ì �� (Ì �� '�L �� '�L ��      >    , � � �� � ��  8 �  8 � �      >    , $d L �0 L �0 ( $d ( $d L      >    , 
�� � �� � �� �� 
�� �� 
�� �      >    , v� a| �� a| �� m4 v� m4 v� a|      >    , '�@   ('L   ('L � '�@ � '�@        >    , � #�� <� #�� <� #�| � #�| � #��      >    , ݈ 	�x 	h 	�x 	h 	�0 ݈ 	�0 ݈ 	�x      >    , _� �L l �L l � _� � _� �L      >    , i� � � � � �� i� �� i� �      >    , �4 � �  � �  �� �4 �� �4 �      >    , ��  �� L  �� L  �8 ��  �8 ��  ��      >    , �< ��  � ��  � �� �< �� �< ��      >    , )� �8 X� �8 X� � )� � )� �8      >    , !?� #�� "Ep #�� "Ep #� !?� #� !?� #��      >    , �X Z� �� Z� �� fd �X fd �X Z�      >    , -|�  h .,P  h .,P   -|�   -|�  h      >    , '!� 	Ӡ *w 	Ӡ *w 	�X '!� 	�X '!� 	Ӡ      >    , #K( >4 %
l >4 %
l I� #K( I� #K( >4      >    , h   ׬   ׬ � h � h        >    , �L `< � `< � k� �L k� �L `<      >    , s� Ҥ �8 Ҥ �8 �\ s� �\ s� Ҥ      >    , �� �8 h �8 h � �� � �� �8      >    , �| �l �x �l �x �$ �| �$ �| �l      >    , �� !Kp 	`d !Kp 	`d !W( �� !W( �� !Kp      >    , $� %�\  %�\  %� $� %� $� %�\      >    , E� � "p � "p �� E� �� E� �      >    ,  | � �p � �p ��  | ��  | �      >    , =� d� �L d� �L p� =� p� =� d�      >    , '�p  � (��  � (��  �H '�p  �H '�p  �      >    , P � J0 � J0 �� P �� P �      >    , >x 0� u( 0� u( <d >x <d >x 0�      >    , ,4 � ,v� � ,v� < ,4 < ,4 �      >    , %` ȼ %}� ȼ %}� �t %` �t %` ȼ      >    , �8 &'� kd &'� kd &3L �8 &3L �8 &'�      >    , �P !�( '� !�( '� !�� �P !�� �P !�(      >    , }  	� �� 	� �� X }  X }  	�      >    , Lp �� � �� � �H Lp �H Lp ��      >    , 
� v� X( v� X( �� 
� �� 
� v�      >    , �� %�L �d %�L �d %� �� %� �� %�L      >    , (� �T �t �T �t � (� � (� �T      >    , �X %�\ l %�\ l %� �X %� �X %�\      >    , N@ @p U� @p U� L( N@ L( N@ @p      >    , 
T� �� %� �� %� �t 
T� �t 
T� ��      >    , +| 28 +�� 28 +�� =� +| =� +| 28      >    ,  � �� � �� ��  ��  �      >    , (X  � (�  � (�  �� (X  �� (X  �      >    , (�� #�� +|� #�� +|� #�| (�� #�| (�� #��      >    , �� i� - i� - u� �� u� �� i�      >    , �  @p � @p � L( �  L( �  @p      >    , "7� �h %� �h %� �  "7� �  "7� �h      >    , y4 i� �� i� �� u� y4 u� y4 i�      >    , 
� =� 8 =� 8 I� 
� I� 
� =�      >    , )�   *�   *� � )� � )�        >    , !T  � S�  � S�  �H !T  �H !T  �      >    , �� b� �� b� �� nX �� nX �� b�      >    , =� i� d� i� d� u� =� u� =� i�      >    ,  �t 	� !.$ 	� !.$ �  �t �  �t 	�      >    , M  %�\ �4 %�\ �4 %� M  %� M  %�\      >    , �� d� �� d� �� p� �� p� �� d�      >    , �4 �, � �, � �� �4 �� �4 �,      >    , (�p ;� )) ;� )) GH (�p GH (�p ;�      >    ,  �< � !� � !� ��  �< ��  �< �      >    , 	'�  d 
f  d 
f  	'�  	'�  d      >    , &� <h (Z <h (Z H  &� H  &� <h      >    , "�4 r� "� r� "� ~d "�4 ~d "�4 r�      >    , 	�l T@ 	�� T@ 	�� _� 	�l _� 	�l T@      >    , �� eD �x eD �x p� �� p� �� eD      >    , %!� >4 &)� >4 &)� I� %!� I� %!� >4      >    , �\ �T 	V� �T 	V� � �\ � �\ �T      >    , ,$� $ -$� $ -$� "� ,$� "� ,$� $      >    , !�p x "U x "U '0 !�p '0 !�p x      >    ,  t� 
ш  �x 
ш  �x 
�@  t� 
�@  t� 
ш      >    , ֈ ٜ $� ٜ $� �T ֈ �T ֈ ٜ      >    , �\ 	f@ _  	f@ _  	q� �\ 	q� �\ 	f@      >    , dH ;� � ;� � GH dH GH dH ;�      >    , { 	�� ,X 	�� ,X 
� { 
� { 	��      >    , _D 
= � 
= � 
H� _D 
H� _D 
=      >    , ,| JT ,�( JT ,�( V ,| V ,| JT      >    , ( ed t4 ed t4 q ( q ( ed      >    , *�@ �\ +�� �\ +�� � *�@ � *�@ �\      >    , P4 �� � �� � �D P4 �D P4 ��      >    , �X �  �  �@ �X �@ �X �      >    , R  � �h  � �h  �H R  �H R  �      >    , )�D � )�$ � )�$ �� )�D �� )�D �      >    , #d� #�� #� #�� #� #� #d� #� #d� #��      >    , !~8   "�   "� � !~8 � !~8        >    , y %�\ &� %�\ &� %� y %� y %�\      >    , �X � +8 � +8 �� �X �� �X �      >    , ?� �� �� �� �� �| ?� �| ?� ��      >    , )�� �� *L �� *L �� )�� �� )�� ��      >    ,  � !� #ݤ !� #ݤ !��  � !��  � !�      >    , � %$ �� %$ �� %!� � %!� � %$      >    , $�X a| %5d a| %5d m4 $�X m4 $�X a|      >    , � O �< O �< Z� � Z� � O      >    , -�l #� . #� . /H -�l /H -�l #�      >    , �D !�L �� !�L �� !� �D !� �D !�L      >    , + !�\ { !�\ { " + " + !�\      >    , q   � �H  � �H d q  d q   �      >    , +< 4 g� 4 g� ?� +< ?� +< 4      >    , }h z� $ z� $ �X }h �X }h z�      >    , �X �� `� �� `� �� �X �� �X ��      >    , �( 
��  Sd 
��  Sd 
�H �( 
�H �( 
��      >    , L� � Ѩ � Ѩ � L� � L� �      >    , � �� A� �� A� �� � �� � ��      >    , 5� s �� s �� ~� 5� ~� 5� s      >    , �8 �� �( �� �( �| �8 �| �8 ��      >    , � i, GD i, GD t� � t� � i,      >    , �< 	?0 	� 	?0 	� 	J� �< 	J� �< 	?0      >    , � � d � d �� � �� � �      >    , )� 	�P +Y� 	�P +Y� 	� )� 	� )� 	�P      >    , � � �  � �  $d � $d � �      >    , d� �D dH �D dH �� d� �� d� �D      >    , �� �� cp �� cp �� �� �� �� ��      >    , ,�D   -G�   -G� � ,�D � ,�D        >    , t�  d ��  d ��  t�  t�  d      >    , &H� �� 'k� �� 'k� �| &H� �| &H� ��      >    , (-( � (� � (� �� (-( �� (-( �      >    , i !�L  � !�L  � !� i !� i !�L      >    , $�p a� &l a� &l m� $�p m� $�p a�      >    , .� $  ._ $  ._ $+� .� $+� .� $       >    , [� �� _� �� _� �| [� �| [� ��      >    , )�T  �� *ڴ  �� *ڴ  �8 )�T  �8 )�T  ��      >    , !� �h "� �h "� �  !� �  !� �h      >    , +� 
d( 	� 
d( 	� 
o� +� 
o� +� 
d(      >    , �� �� �� �� �� �� �� �� �� ��      >    , s� �( �$ �( �$ �� s� �� s� �(      >    , 
j ~@ �� ~@ �� �� 
j �� 
j ~@      >    , v� Z� �� Z� �� fd v� fd v� Z�      >    , �@ &l � &l � &$ �@ &$ �@ &l      >    , �p � ,8 � ,8 �� �p �� �p �      >    , tX �� � �� � �T tX �T tX ��      >    , S� � �H � �H �@ S� �@ S� �      >    , ]� 	� ~� 	� ~� X ]� X ]� 	�      >    , �0 \ �$ \ �$   �0   �0 \      >    , �� 	�P �| 	�P �| 	� �� 	� �� 	�P      >    , +�H � -� � -� �X +�H �X +�H �      >    , ,�� � -�� � -��  8 ,��  8 ,�� �      >    , 4p �� �, �� �, �| 4p �| 4p ��      >    , 
L %�\ #� %�\ #� %� 
L %� 
L %�\      >    , $=X #�� %H #�� %H #�| $=X #�| $=X #��      >    , �h $ Ƥ $ Ƥ "� �h "� �h $      >    , ߠ 	f@ 
F� 	f@ 
F� 	q� ߠ 	q� ߠ 	f@      >    , � >4 <� >4 <� I� � I� � >4      >    , "�� �\ #� �\ #� � "�� � "�� �\      >    , !�@ `< !�  `< !�  k� !�@ k� !�@ `<      >    ,  �D b�  �$ b�  �$ nX  �D nX  �D b�      >    , �� ø � ø � �p �� �p �� ø      >    , �` �4 @ �4 @ �� �` �� �` �4      >    , #�� 	�P %�X 	�P %�X 	� #�� 	� #�� 	�P      >    , )� �� *�@ �� *�@ �T )� �T )� ��      >    , E� eD C� eD C� p� E� p� E� eD      >    , +�p |� ,�� |� ,�� �D +�p �D +�p |�      >    , $� !�< %�$ !�< %�$ !�� $� !�� $� !�<      >    , !�l �T !�@ �T !�@ � !�l � !�l �T      >    , ې `� �� `� �� l� ې l� ې `�      >    , Vx �T � �T � � Vx � Vx �T      >    , !�H ~� ".  ~� ".  �� !�H �� !�H ~�      >    , $� �� $�� �� $�� �L $� �L $� ��      >    , &^D �� ' �� ' �T &^D �T &^D ��      >    , )  	?0 *B\ 	?0 *B\ 	J� )  	J� )  	?0      >    , 	�� |( � |( � �� 	�� �� 	�� |(      >    , �� �� �| �� �| �� �� �� �� ��      >    , �� 	f@ �  	f@ �  	q� �� 	q� �� 	f@      >    , & [ T� [ T� f� & f� & [      >    , 	{� �d 
D �d 
D � 	{� � 	{� �d      >    , � &l 7� &l 7� &$ � &$ � &l      >    , Z� ,� �� ,� �� 8� Z� 8� Z� ,�      >    , 	�h �� � �� � ̨ 	�h ̨ 	�h ��      >    , 	 � 7� � 7� �� 	 �� 	 �      >    , $E( �8 %�( �8 %�( � $E( � $E( �8      >    , (� B�  � B�  � N@ (� N@ (� B�      >    , 9, w  �� w  �� �� 9, �� 9, w       >    , (T8 >4 )� >4 )� I� (T8 I� (T8 >4      >    , $� �4 $�  �4 $�  �� $� �� $� �4      >    , "3� ;� $ � ;� $ � GH "3� GH "3� ;�      >    , 1< �D �  �D �  �� 1< �� 1< �D      >    , �x 4 �0 4 �0 ?� �x ?� �x 4      >    , (� �L W� �L W� � (� � (� �L      >    , z� 	f@ � 	f@ � 	q� z� 	q� z� 	f@      >    , �( >4 u� >4 u� I� �( I� �( >4      >    , (� �d )+ �d )+ � (� � (� �d      >    , $�� �l &x �l &x �$ $�� �$ $�� �l      >    , �P H ~@ H ~@ )  �P )  �P H      >    , - ʬ -A� ʬ -A� �d - �d - ʬ      >    , ,|� �( -Ux �( -Ux �� ,|� �� ,|� �(      >    , &i� �� &�� �� &�� � &i� � &i� ��      >    , =� 1 
� 1 
� <� =� <� =� 1      >    , ʰ i� �P i� �P u� ʰ u� ʰ i�      >    , � 	?0 X� 	?0 X� 	J� � 	J� � 	?0      >    , �� �  �� �  �� �� �� �� �� �       >    , -�D J� -�� J� -�� VX -�D VX -�D J�      >    , dH :l �  :l �  F$ dH F$ dH :l      >    , ,\ 	?0 � 	?0 � 	J� ,\ 	J� ,\ 	?0      >    , �4 	�� �$ 	�� �$ 
� �4 
� �4 	��      >    , 
 r� 4� r� 4� ~d 
 ~d 
 r�      >    , -� !�\ }� !�\ }� " -� " -� !�\      >    , %< �4 �$ �4 �$ �� %< �� %< �4      >    , �� �� !�  �� !�  �� �� �� �� ��      >    , 5� �T M  �T M  � 5� � 5� �T      >    , �` ', @ ', @ 2� �` 2� �` ',      >    , 	X �� 88 �� 88 �� 	X �� 	X ��      >    , AD �4 �d �4 �d �� AD �� AD �4      >    , "�� �� #�x �� #�x �T "�� �T "�� ��      >    ,  � $  %�  $  %�  $+�  � $+�  � $       >    , )� � +d � +d < )� < )� �      >    , *��  d +��  d +��  *��  *��  d      >    , �   �h   �h � � � �        >    , X� %$ �� %$ �� %!� X� %!� X� %$      >    , �� �� �d �� �d l �� l �� ��      >    , �� eD  � eD  � p� �� p� �� eD      >    , *�� �� +� �� +� �� *�� �� *�� ��      >    , �� 	׈ Ը 	׈ Ը 	�@ �� 	�@ �� 	׈      >    , (� !x "�0 !x "�0 -0 (� -0 (� !x      >    , \4 � +� � +� +� \4 +� \4 �      >    , �d � 'T � 'T � �d � �d �      >    , 3� �| fd �| fd �4 3� �4 3� �|      >    , � �h �� �h �� �  � �  � �h      >    , h �� !� �� !� �� h �� h ��      >    , �� %�\ `` %�\ `` %� �� %� �� %�\      >    , �� �� �� �� �� �D �� �D �� ��      >    , ,�� �� -l� �� -l� �T ,�� �T ,�� ��      >    , &F� :l &w� :l &w� F$ &F� F$ &F� :l      >    , y4 #� I� #� I� /D y4 /D y4 #�      >    , �(   ��   �� � �( � �(        >    , vp �� x@ �� x@ � vp � vp ��      >    , � ', ( ', ( 2� � 2� � ',      >    , R( #�� � #�� � #� R( #� R( #��      >    , 	/� "� 	�� "� 	�� "�� 	/� "�� 	/� "�      >    , �X !�L t� !�L t� !� �X !� �X !�L      >    , +o$ � ,B � ,B � +o$ � +o$ �      >    ,  �� �� !�� �� !�� �|  �� �|  �� ��      >    , *�P b� +�d b� +�d nX *�P nX *�P b�      >    , +�� [ +�  [ +�  f� +�� f� +�� [      >    , +_� !�L ,g0 !�L ,g0 !� +_� !� +_� !�L      >    , iL d� � d� � p� iL p� iL d�      >    , �P ( �x ( �x � �P � �P (      >    , 
B� 4 
�� 4 
�� ?� 
B� ?� 
B� 4      >    , $�� �� $ی �� $ی �| $�� �| $�� ��      >    , �, ( �� ( �� � �, � �, (      >    , )!L ;� *!( ;� *!( GH )!L GH )!L ;�      >    , �h f< g\ f< g\ q� �h q� �h f<      >    , ^  ;� �@ ;� �@ GH ^  GH ^  ;�      >    , �� �l e  �l e  �$ �� �$ �� �l      >    ,  �< 	׈ & � 	׈ & � 	�@  �< 	�@  �< 	׈      >    , )l �� � �� � �� )l �� )l ��      >    , '� �� '�@ �� '�@ �� '� �� '� ��      >    , 	�� J� 	�d J� 	�d VT 	�� VT 	�� J�      >    ,  :  #��  � #��  � #�  :  #�  :  #��      >    , +� �� 	�p �� 	�p �t +� �t +� ��      >    , � �� �  �� �  �� � �� � ��      >    , ?t eD d eD d p� ?t p� ?t eD      >    , dp >4 	  >4 	  I� dp I� dp >4      >    , �� �� �  �� �  �� �� �� �� ��      >    , Rp 	� � 	� � X Rp X Rp 	�      >    , �| |� 	 |� 	 �D �| �D �| |�      >    , 
�x ( 
�X ( 
�X � 
�x � 
�x (      >    , /� �� � �� � �T /� �T /� ��      >    , 
1` �� 
h �� 
h �T 
1` �T 
1` ��      >    , l� a| y� a| y� m4 l� m4 l� a|      >    , �� �( 4� �( 4� �� �� �� �� �(      >    , �T !�\ �� !�\ �� " �T " �T !�\      >    , #� #�� #M #�� #M #� #� #� #� #��      >    , �� ', ;h ', ;h 2� �� 2� �� ',      >    , �� 
�h �H 
�h �H 
�  �� 
�  �� 
�h      >    , 4p �$ �� �$ �� �� 4p �� 4p �$      >    , �� 	� 80 	� 80 X �� X �� 	�      >    , 	bX \ 
5H \ 
5H  	bX  	bX \      >    , �P |� �  |� �  �D �P �D �P |�      >    , �\ 	f@ iL 	f@ iL 	q� �\ 	q� �\ 	f@      >    , � �� � �� � �� � �� � ��      >    , � �� <� �� <� 	 � � 	 � � ��      >    , 1� �x �� �x �� �0 1� �0 1� �x      >    , � F� \ F� \ Rp � Rp � F�      >    , 	� �� � �� � � 	� � 	� ��      >    , ]0 ٜ � ٜ � �T ]0 �T ]0 ٜ      >    , � �� �x �� �x �x � �x � ��      >    ,  "�� � "�� � "��  "��  "��      >    , (�X �T )H\ �T )H\ � (�X � (�X �T      >    , #�� �� '�� �� '�� �� #�� �� #�� ��      >    , �  �� ��  �� ��  Ơ �  Ơ �  ��      >    , � :l �� :l �� F$ � F$ � :l      >    , #7� Đ $٘ Đ $٘ �H #7� �H #7� Đ      >    , T  � h  � h  �H T  �H T  �      >    , O< \ �� \ ��   O<   O< \      >    , � � 	�h � 	�h  8 �  8 � �      >    , '� j� (� j� (� vp '� vp '� j�      >    , �� 	j( ݨ 	j( ݨ 	u� �� 	u� �� 	j(      >    , T` v� �� v� �� �� T` �� T` v�      >    , V4  d Bd  d Bd  V4  V4  d      >    , �0 "�D �8 "�D �8 "�� �0 "�� �0 "�D      >    , �� /� �� /� �� ;� �� ;� �� /�      >    , � 	?0 ,� 	?0 ,� 	J� � 	J� � 	?0      >    , 'P  �� �  �� �  �8 'P  �8 'P  ��      >    , , 84 8 84 8 C� , C� , 84      >    , 4P �4 i �4 i �� 4P �� 4P �4      >    , *�� :l +�@ :l +�@ F$ *�� F$ *�� :l      >    , 'e� � (�� � (�� �� 'e� �� 'e� �      >    , � ��  :  ��  :  �� � �� � ��      >    , 5� � V� � V� �� 5� �� 5� �      >    , 1� #�� E, #�� E, #� 1� #� 1� #��      >    , �X O  P O  P Z� �X Z� �X O      >    , H� �� �� �� �� �T H� �T H� ��      >    , h �� �� �� �� �| h �| h ��      >    , #�� �� &d  �� &d  �� #�� �� #�� ��      >    , �� %�\ W %�\ W %� �� %� �� %�\      >    , "� �D #EL �D #EL �� "� �� "� �D      >    , 2\ #� А #� А /� 2\ /� 2\ #�      >    , *ܨ �� +� �� +� �T *ܨ �T *ܨ ��      >    ,  � � � � ��  ��  �      >    , � � �� � ��  8 �  8 � �      >    , � O � O � Z� � Z� � O      >    , 6< 	� !� 	� !� X 6< X 6< 	�      >    , #�0  � #�  � #�  �H #�0  �H #�0  �      >    , y� �� �p �� �p �| y� �| y� ��      >    , #�� 	?0 %F� 	?0 %F� 	J� #�� 	J� #�� 	?0      >    , #�0 \ $�4 \ $�4  #�0  #�0 \      >    , �� :l tT :l tT F$ �� F$ �� :l      >    , &i� JT *�@ JT *�@ V &i� V &i� JT      >    , � , �� , ��  � �  � � ,      >    , $�h #�� %�� #�� %�� #� $�h #� $�h #��      >    , "p �| =� �| =� 4 "p 4 "p �|      >    , ��   ��   �� � �� � ��        >    , !� H #+� H #+� )  !� )  !� H      >    , �� �@ �$ �@ �$ �� �� �� �� �@      >    ,  	�P A� 	�P A� 	�  	�  	�P      >    , *�� �� *�` �� *�` �| *�� �| *�� ��      >    , -�D �� .A� �� .A� �T -�D �T -�D ��      >    , < \ O� \ O�  <  < \      >    , )�p ', +@ ', +@ 2� )�p 2� )�p ',      >    , �� #�� {L #�� {L #� �� #� �� #��      >    , �|   ��   �� � �| � �|        >    , $7| � %0 � %0 �� $7| �� $7| �      >    , `` �T �  �T �  � `` � `` �T      >    , )� �� )� �� )� �T )� �T )� ��      >    , )| ?t )�( ?t )�( K, )| K, )| ?t      >    , �� �8 _@ �8 _@ � �� � �� �8      >    , !� [ "�� [ "�� f� !� f� !� [      >    , ��  � �(  � �(  �H ��  �H ��  �      >    , �� :l �p :l �p F$ �� F$ �� :l      >    , -Ux :l .�P :l .�P F$ -Ux F$ -Ux :l      >    , �@ :l �� :l �� F$ �@ F$ �@ :l      >    , +�, �8 ,�` �8 ,�` � +�, � +�, �8      >    , eh �� �� �� �� �T eh �T eh ��      >    , � #�� �  #�� �  #� � #� � #��      >    , tX � GH � GH �� tX �� tX �      >    , 
B� &l s� &l s� &$ 
B� &$ 
B� &l      >    , �� #�� � #�� � #� �� #� �� #��      >    , � %�$ � %�$ � %�� � %�� � %�$      >    , �   �0   �0 � � � �        >    , � %�\ �� %�\ �� %� � %� � %�\      >    , %�` �� %�@ �� %�@ �� %�` �� %�` ��      >    , #�� �� $� �� $� �T #�� �T #�� ��      >    , �   U�   U� � � � �        >    , *�P � -K� � -K� �� *�P �� *�P �      >    , �$ &l o &l o &$ �$ &$ �$ &l      >    , 	?0 %o� � %o� � %{� 	?0 %{� 	?0 %o�      >    , �, �� /� �� /� �� �, �� �, ��      >    , C8 � � � � �� C8 �� C8 �      >    , �, �� �� �� �� �� �, �� �, ��      >    , ��  �` ��  �` ��  � ��  � ��  �`      >    , �, \ !	 \ !	   �,   �, \      >    , < $f\ 0 $f\ 0 $r < $r < $f\      >    , �| $��  �� $��  �� $�< �| $�< �| $��      >    , 7� d�  � d�  � pl 7� pl 7� d�      >    , '� �$ '�D �$ '�D �� '� �� '� �$      >    , % � :l &� :l &� F$ % � F$ % � :l      >    , Y� �4 �� �4 �� �� Y� �� Y� �4      >    , � "� �H "� �H "$< � "$< � "�      >    , ,\ #�� �x #�� �x #� ,\ #� ,\ #��      >    , (�<  d *~�  d *~�  (�<  (�<  d      >    , !� %�\ !�, %�\ !�, %� !� %� !� %�\      >    , **� = *�� = *�� H� **� H� **� =      >    , $`� `< %j  `< %j  k� $`� k� $`� `<      >    , Fp � _� � _� �� Fp �� Fp �      >    , U| �  � �  � �� U| �� U| �      >    , �P 	� ( 	� ( X �P X �P 	�      >    , �P [ �x [ �x f� �P f� �P [      >    , l� S� � S� � _� l� _� l� S�      >    , %w� ;� &� ;� &� GH %w� GH %w� ;�      >    , {t �� , �� , �D {t �D {t ��      >    ,  � @p � @p � L(  � L(  � @p      >    , vp H � H � )  vp )  vp H      >    , )� �� +O� �� +O� �� )� �� )� ��      >    , E�  � ��  � ��  �H E�  �H E�  �      >    , l�  � .P  � .P  �H l�  �H l�  �      >    , N� z� �( z� �( �X N� �X N� z�      >    , �X 	�P rd 	�P rd 	� �X 	� �X 	�P      >    , �T 4 �� 4 �� ?� �T ?� �T 4      >    , � \ =� \ =�   �   � \      >    , H #�� @( #�� @( #� H #� H #��      >    , � !�< #$ !�< #$ !�� � !�� � !�<      >    , ,Ш 	f@ -� 	f@ -� 	q� ,Ш 	q� ,Ш 	f@      >    , *�\ � ,4h � ,4h �� *�\ �� *�\ �      >    , �� �, �H �, �H �� �� �� �� �,      >    , �4 $  � $  � $+� �4 $+� �4 $       >    , h � �d � �d &| h &| h �      >    , "� � #�� � #�� �� "� �� "� �      >    , Fl ;� �| ;� �| G� Fl G� Fl ;�      >    , ڸ   .�   .� � ڸ � ڸ        >    , �� �D ̀ �D ̀ �� �� �� �� �D      >    , �� #l  �� #l  �� #"$ �� #"$ �� #l      >    , �P ٜ ]T ٜ ]T �T �P �T �P ٜ      >    , �p %�L ! %�L ! %� �p %� �p %�L      >    , "?� `< "nt `< "nt k� "?� k� "?� `<      >    , \� &l �\ &l �\ &$ \� &$ \� &l      >    , '< � 'J� � 'J� �� '< �� '< �      >    , ��   �   � � �� � ��        >    , E� #�� "�� #�� "�� #�T E� #�T E� #��      >    ,  ?�  � !��  � !��  �H  ?�  �H  ?�  �      >    , �� :l <� :l <� F$ �� F$ �� :l      >    , μ !�L �� !�L �� !� μ !� μ !�L      >    , 	\| !�\ 
� !�\ 
� " 	\| " 	\| !�\      >    , �0 �� � �� � �T �0 �T �0 ��      >    , a �� � �� � �� a �� a ��      >    , �� � 	n � 	n %� �� %� �� �      >    , �X b� � b� � nX �X nX �X b�      >    , *@ �4 Y  �4 Y  �� *@ �� *@ �4      >    , �   �   � � � � �        >    , �d �� �$ �� �$ � �d � �d ��      >    , ( < h (�8 h (�8   ( <   ( < h      >    , �� !8 #�  !8 #�  !� �� !� �� !8      >    , �@ 	��  	��  	׈ �@ 	׈ �@ 	��      >    , 	j( � 	�� � 	�� +� 	j( +� 	j( �      >    , �l #�� 0 #�� 0 #�| �l #�| �l #��      >    , )mx $G .j� $G .j� $R� )mx $R� )mx $G      >    , �` �� �@ �� �@ �@ �` �@ �` ��      >    , �� d� ˨ d� ˨ pl �� pl �� d�      >    , )�� �$ *Y� �$ *Y� �� )�� �� )�� �$      >    , �P 
� � 
� � 
%� �P 
%� �P 
�      >    , � � �\ � �\ �� � �� � �      >    , �� �� e@ �� e@ �l �� �l �� ��      >    , 7� 	�` XH 	�` XH 	� 7� 	� 7� 	�`      >    , $�| "�� &$ "�� &$ "�� $�| "�� $�| "��      >    , "�x !�< "�@ !�< "�@ !�� "�x !�� "�x !�<      >    , 	� �� e@ �� e@ �� 	� �� 	� ��      >    , "�  � #��  � #��  �H "�  �H "�  �      >    , +�� �4 ,�� �4 ,�� � +�� � +�� �4      >    , /h �T ^H �T ^H � /h � /h �T      >    , !b� x !�  x !�  '0 !b� '0 !b� x      >    , �� eD  4$ eD  4$ p� �� p� �� eD      >    , | F� �� F� �� Rl | Rl | F�      >    , �h %�\ a� %�\ a� %� �h %� �h %�\      >    , �l Ҥ �( Ҥ �( �\ �l �\ �l Ҥ      >    , 
�< !�, d !�, d !�� 
�< !�� 
�< !�,      >    , .P a| �� a| �� m4 .P m4 .P a|      >    , �0 p$ �  p$ �  {� �0 {� �0 p$      >    , �< \ �� \ ��  �<  �< \      >    , �� !�T �8 !�T �8 !� �� !� �� !�T      >    ,  ¸ �� "� �� "� �T  ¸ �T  ¸ ��      >    , �� �l 	� �l 	� �$ �� �$ �� �l      >    , '�( �� (PP �� (PP �| '�( �| '�( ��      >    , '14 	� '�� 	� '�� x '14 x '14 	�      >    , $�H �T %H �T %H � $�H � $�H �T      >    , 6  �| ̄ �| ̄ �4 6  �4 6  �|      >    , �� %�\ �� %�\ �� %� �� %� �� %�\      >    , > [| �� [| �� g4 > g4 > [|      >    , &�P �l '0 �l '0 �$ &�P �$ &�P �l      >    , !� �� %5d �� %5d | !� | !� ��      >    , 
h e� 
ϔ e� 
ϔ q� 
h q� 
h e�      >    , � �� 5  �� 5  ݈ � ݈ � ��      >    , �8 �8  �8  � �8 � �8 �8      >    , "�p #�� $?L #�� $?L #�| "�p #�| "�p #��      >    , /� =� pL =� pL I� /� I� /� =�      >    , 0� Đ ed Đ ed �H 0� �H 0� Đ      >    , �� 0� �� 0� �� <h �� <h �� 0�      >    , �� $ �\ $ �\ "� �� "� �� $      >    , )�� �� *�� �� *�� �D )�� �D )�� ��      >    , %l   '��   '�� � %l � %l        >    , �� [ �� [ �� f� �� f� �� [      >    , C� � �� � ��  8 C�  8 C� �      >    , �� $�� L� $�� L� $�< �� $�< �� $��      >    , �4 �� � �� � �l �4 �l �4 ��      >    , &4 "�� �\ "�� �\ "�� &4 "�� &4 "��      >    , � �d  M� �d  M� � � � � �d      >    , '3( 
( (�� 
( (�� � '3( � '3( 
(      >    , ,d �@ ,:D �@ ,:D �� ,d �� ,d �@      >    , �  ި �  ި �  �` �  �` �  ި      >    , r� �� � �� � �| r� �| r� ��      >    , ƀ ~� �` ~� �` �\ ƀ �\ ƀ ~�      >    , �P "� �, "� �, "$< �P "$< �P "�      >    , �@ ( d ( d � �@ � �@ (      >    , j� � l� � l� �� j� �� j� �      >    , h� 	� �� 	� �� X h� X h� 	�      >    , �� �8 � �8 � � �� � �� �8      >    , eH � k  � k  �� eH �� eH �      >    , /D 4 � 4 � ?� /D ?� /D 4      >    , SH �( S$ �( S$ �� SH �� SH �(      >    , < �� r� �� r� �t < �t < ��      >    , 
  � T@ � T@ &| 
  &| 
  �      >    , � � 	�  � 	�  �� � �� � �      >    , � %�\ �� %�\ �� %� � %� � %�\      >    , 
�� 
= Rp 
= Rp 
H� 
�� 
H� 
�� 
=      >    , 
 %�$ 
s� %�$ 
s� %�� 
 %�� 
 %�$      >    , 4 %�\ �P %�\ �P %� 4 %� 4 %�\      >    , 	�< |� �\ |� �\ �D 	�< �D 	�< |�      >    , � !�, 	�P !�, 	�P !�� � !�� � !�,      >    , +֨ �� ,�x �� ,�x �T +֨ �T +֨ ��      >    , $�@ L %x L %x W� $�@ W� $�@ L      >    , ׄ �� �0 �� �0 �T ׄ �T ׄ ��      >    , �� #�� �� #�� �� #� �� #� �� #��      >    , r� !�L Q� !�L Q� !� r� !� r� !�L      >    , i0 �( �, �( �, �� i0 �� i0 �(      >    , �� ( =� ( =� � �� � �� (      >    , 6� %�\ � %�\ � %� 6� %� 6� %�\      >    , +cl i� ,<8 i� ,<8 u� +cl u� +cl i�      >    , � �  7� �  7� �� � �� � �       >    , �  :l � :l � F$ �  F$ �  :l      >    , � !8 �$ !8 �$ !� � !� � !8      >    , �, !�< � !�< � !�� �, !�� �, !�<      >    ,  zt %�L !f� %�L !f� %�  zt %�  zt %�L      >    , �D "� '� "� '� "�� �D "�� �D "�      >    , F� d� �� d� �� p� F� p� F� d�      >    , +�� 	p ,� 	p ,� 	{� +�� 	{� +�� 	p      >    , ?x %�\ �  %�\ �  %� ?x %� ?x %�\      >    , )6� �0 )e� �0 )e� �� )6� �� )6� �0      >    , &Ǽ 
� (�$ 
� (�$ 
+� &Ǽ 
+� &Ǽ 
�      >    , "Z� 
� $T� 
� $T� � "Z� � "Z� 
�      >    , q  � &�  � &�  �H q  �H q  �      >    , �@ �� �� �� �� �� �@ �� �@ ��      >    , ��  d �  d �  ��  ��  d      >    , 
�� d� Ǡ d� Ǡ pl 
�� pl 
�� d�      >    , "�P �4 #�( �4 #�( �� "�P �� "�P �4      >    ,   � c( � c( �   �   �      >    , �p [| �P [| �P g4 �p g4 �p [|      >    , � 	f@ �� 	f@ �� 	q� � 	q� � 	f@      >    , *c� !�< +�L !�< +�L !�� *c� !�� *c� !�<      >    , � �� T� �� T� �� � �� � ��      >    , �� �� � �� � �� �� �� �� ��      >    , wh 	Ӡ iP 	Ӡ iP 	�X wh 	�X wh 	Ӡ      >    , #^� H $%� H $%� )  #^� )  #^� H      >    , �� i� "� i� "� u� �� u� �� i�      >    , < %�\ � %�\ � %� < %� < %�\      >    , h �� :l �� :l �| h �| h ��      >    , '�� ?t (� ?t (� K, '�� K, '�� ?t      >    , g  �� vp  �� vp  Ơ g  Ơ g  ��      >    , =� m� � m� � y| =� y| =� m�      >    , _H 4 e  4 e  ?� _H ?� _H 4      >    , m �� Ҥ �� Ҥ �� m �� m ��      >    ,   � �  � �  �H   �H   �      >    , 4 � �� � �� �� 4 �� 4 �      >    , 	4 � � � � � 	4 � 	4 �      >    , � 4 fd 4 fd ?� � ?� � 4      >    , /H  � 3  � 3  �H /H  �H /H  �      >    , � �� > �� > �� � �� � ��      >    , 	��  � 
^L  � 
^L  �H 	��  �H 	��  �      >    , �T d� ] d� ] p� �T p� �T d�      >    , �( :l �� :l �� F$ �( F$ �( :l      >    , 	3x d� 	�� d� 	�� p� 	3x p� 	3x d�      >    , � �$ 5h �$ 5h �� � �� � �$      >    , <� � �L � �L �� <� �� <� �      >    , ,�� �8 -�L �8 -�L � ,�� � ,�� �8      >    , ,�@ >4 -ΐ >4 -ΐ I� ,�@ I� ,�@ >4      >    , ٜ !�< %� !�< %� !�� ٜ !�� ٜ !�<      >    ,  �$ D0  � D0  � O�  �$ O�  �$ D0      >    , � �8 2� �8 2� � � � � �8      >    , ' H � H � )  ' )  ' H      >    , @ , ` , `  � @  � @ ,      >    , � 	f@ �, 	f@ �, 	q� � 	q� � 	f@      >    , #�� ( %^h ( %^h � #�� � #�� (      >    , (�� �� )�� �� )�� �D (�� �D (�� ��      >    , gX %�\ �� %�\ �� %� gX %� gX %�\      >    , %/� =� %Ә =� %Ә I� %/� I� %/� =�      >    , r� � � � �  8 r�  8 r� �      >    , b !� � !� � !�� b !�� b !�      >    , �( 	f@ ~� 	f@ ~� 	q� �( 	q� �( 	f@      >    , �� !�L �� !�L �� !� �� !� �� !�L      >    ,  �  "�D #l\ "�D #l\ "��  �  "��  �  "�D      >    , � �� �� �� �� �T � �T � ��      >    , )R  �� +2� �� +2� �p )R  �p )R  ��      >    , 
� S� ,4 S� ,4 _� 
� _� 
� S�      >    , 	{�  �� 
�H  �� 
�H  �8 	{�  �8 	{�  ��      >    , ]� =� 0� =� 0� I� ]� I� ]� =�      >    , -�P d� .S` d� .S` pl -�P pl -�P d�      >    , P 't x 't x 3, P 3, P 't      >    , @�   ɔ   ɔ � @� � @�        >    , � �� ְ �� ְ ߜ � ߜ � ��      >    , &ɰ !�\ (:� !�\ (:� " &ɰ " &ɰ !�\      >    , nX =� AH =� AH I� nX I� nX =�      >    , '��  N  (
   N  (
   Y� '��  Y� '��  N       >    ,  �8 �x �8 �x �  �  �8      >    , +�` ', ,�  ', ,�  2� +�` 2� +�` ',      >    , C�   �L   �L � C� � C�        >    , j� !� �D !� �D !�� j� !�� j� !�      >    , �0 %�L �d %�L �d %� �0 %� �0 %�L      >    , Đ � (, � (, 	� Đ 	� Đ �      >    , � #�� 	� #�� 	� #�| � #�| � #��      >    , "Ep |� #^� |� #^� �D "Ep �D "Ep |�      >    , 
�� 	?0 \ 	?0 \ 	J� 
�� 	J� 
�� 	?0      >    , �,  �� �(  �� �(  �8 �,  �8 �,  ��      >    , 	T� �� 	�8 �� 	�8 А 	T� А 	T� ��      >    , @� �� w� �� w� �� @� �� @� ��      >    , rd &l 8 &l 8 &$ rd &$ rd &l      >    , )�� S� *�  S� *�  _� )�� _� )�� S�      >    , "P � 9� � 9� � "P � "P �      >    , +؜ >4 ,S� >4 ,S� I� +؜ I� +؜ >4      >    , ![ �( "�� �( "�� �� ![ �� ![ �(      >    , *�p ;� +�� ;� +�� GH *�p GH *�p ;�      >    , 	�H 6� 
-x 6� 
-x B@ 	�H B@ 	�H 6�      >    , �� �� �H �� �H �� �� �� �� ��      >    , 
� C <� C <� N� 
� N� 
� C      >    , &ɰ � ' ` � ' `  8 &ɰ  8 &ɰ �      >    , !  
A  % � 
A  % � 
L� !  
L� !  
A       >    , &�< "^� (ŀ "^� (ŀ "j� &�< "j� &�< "^�      >    , $� #�� $�L #�� $�L #� $� #� $� #��      >    , �t �( wd �( wd �� �t �� �t �(      >    , 	C �� 	ϸ �� 	ϸ �| 	C �| 	C ��      >    , 	� �� 
� �� 
� �| 	� �| 	� ��      >    , �� �� x �� x �� �� �� �� ��      >    , O� 	f@ 0  	f@ 0  	q� O� 	q� O� 	f@      >    , � �� �@ �� �@ �t � �t � ��      >    , �� �� 	L� �� 	L� �D �� �D �� ��      >    , f� �| �� �| �� 4 f� 4 f� �|      >    , $� �� �$ �� �$ | $� | $� ��      >    , P t� �� t� �� �X P �X P t�      >    , 
�@ !�T  !�T  !� 
�@ !� 
�@ !�T      >    , �� $ �� $ �� "� �� "� �� $      >    , &{� d$ '� d$ '� o� &{� o� &{� d$      >    , B� %�L Z %�L Z %� B� %� B� %�L      >    , �P s �� s �� ~� �P ~� �P s      >    , ̀ !�< \� !�< \� !�� ̀ !�� ̀ !�<      >    , ?t 	�P nT 	�P nT 	� ?t 	� ?t 	�P      >    , +�� `� +� `� +� l� +�� l� +�� `�      >    , ��  �� �  �� �  Ơ ��  Ơ ��  ��      >    , �� 
= �� 
= �� 
H� �� 
H� �� 
=      >    , "7�  � "�  � "�  �H "7�  �H "7�  �      >    , t :l h� :l h� F$ t F$ t :l      >    , h $�� FH $�� FH $�d h $�d h $��      >    , ,@  d -M�  d -M�  ,@  ,@  d      >    , �� � !�� � !�� � �� � �� �      >    , (PP ʬ )g� ʬ )g� �d (PP �d (PP ʬ      >    , ,�� �D ,�� �D ,�� �� ,�� �� ,�� �D      >    , %�p 0� %�P 0� %�P <d %�p <d %�p 0�      >    , - ~@ .08 ~@ .08 �� - �� - ~@      >    , "ph � % � % �� "ph �� "ph �      >    , ,�� �x -�@ �x -�@ �0 ,�� �0 ,�� �x      >    , �� = "�� = "�� H� �� H� �� =      >    , "� a� $�  a� $�  m� "� m� "� a�      >    ,  �| �� '\, �� '\, �L  �| �L  �| ��      >    ,  C� �  r� �  r� ��  C� ��  C� �      >    , ̤ a| C� a| C� m4 ̤ m4 ̤ a|      >    , �d ʬ �� ʬ �� �d �d �d �d ʬ      >    , 4� a| cp a| cp m4 4� m4 4� a|      >    , �p � o� � o� �� �p �� �p �      >    , )y0 �� )�� �� )�� � )y0 � )y0 ��      >    , f� 7� =� 7� =� C< f� C< f� 7�      >    , �� �4 dp �4 dp �� �� �� �� �4      >    , R( �� � �� � �D R( �D R( ��      >    , C� L �� L ��  C�  C� L      >    , �� �� ޤ �� ޤ � �� � �� ��      >    , �� 	Ӡ �� 	Ӡ �� 	�X �� 	�X �� 	Ӡ      >    , 	�� S� 
T� S� 
T� _� 	�� _� 	�� S�      >    ,  �  �� �  �� ø  ø  �       >    , Sh ?t 0 ?t 0 K, Sh K, Sh ?t      >    , �� ( k� ( k� � �� � �� (      >    , ~� �� �� �� �� ̨ ~� ̨ ~� ��      >    , �� "� #EL "� #EL "�� �� "�� �� "�      >    , � $ �� $ �� "� � "� � $      >    , � + �8 + �8 6� � 6� � +      >    , �� 	� �  	� �  X �� X �� 	�      >    , &� �� &�� �� &�� А &� А &� ��      >    , d �� Z� �� Z� �� d �� d ��      >    , 
7< ', s� ', s� 2� 
7< 2� 
7< ',      >    , Ƥ [| �x [| �x g4 Ƥ g4 Ƥ [|      >    , �p �8 �@ �8 �@ � �p � �p �8      >    , �| �� �� �� �� ̨ �| ̨ �| ��      >    , &74  � &��  � &�� � &74 � &74  �      >    , �t �| �� �| �� 4 �t 4 �t �|      >    , 8� #�� :� #�� :� #� 8� #� 8� #��      >    , �  d !r�  d !r�  �  �  d      >    , �� �� >4 �� >4 | �� | �� ��      >    , i0 �� �P �� �P �� i0 �� i0 ��      >    , D @p D� @p D� L( D L( D @p      >    , $E( �$ (o� �$ (o� � $E( � $E( �$      >    , �| �� |( �� |( �T �| �T �| ��      >    , %q� a| &Ǽ a| &Ǽ m4 %q� m4 %q� a|      >    , Q� �� �� �� �� �T Q� �T Q� ��      >    , ۴ "�D AD "�D AD "�� ۴ "�� ۴ "�D      >    , n� �� �h �� �h �� n� �� n� ��      >    , �<  �   �   �H �<  �H �<  �      >    , PX !�L �� !�L �� !� PX !� PX !�L      >    , $'�   $��   $�� � $'� � $'�        >    , '�� $ (yT $ (yT "� '�� "� '�� $      >    , \� � �\ � �\ +� \� +� \� �      >    , D� %�\ �L %�\ �L %� D� %� D� %�\      >    , 'P �D X  �D X  �� 'P �� 'P �D      >    , +�p :l ,�P :l ,�P F$ +�p F$ +�p :l      >    , !�� �� "� �� "� �� !�� �� !�� ��      >    , $0  � &q�  � &q�  � $0  � $0  �      >    , %�� �@ &m� �@ &m� �� %�� �� %�� �@      >    , , �� !�� �� !�� �x , �x , ��      >    , �� �T �� �T �� � �� � �� �T      >    , !�  %�L "� %�L "� %� !�  %� !�  %�L      >    , & #�� &� #�� &� #�| & #�| & #��      >    , �� d� ƀ d� ƀ p� �� p� �� d�      >    , -| �� -�� �� -�� ֬ -| ֬ -| ��      >    , %< [| a� [| a� g4 %< g4 %< [|      >    , "�� ( #�� ( #�� � "�� � "�� (      >    , � #� а #� а /D � /D � #�      >    , .� � �t � �t �� .� �� .� �      >    , k� 	�P �� 	�P �� 	� k� 	� k� 	�P      >    , �, �T � �T � � �, � �, �T      >    , W� � �� � �� �� W� �� W� �      >    , �� �( � �( � �� �� �� �� �(      >    , "�D #� &�d #� &�d /D "�D /D "�D #�      >    , &P� i� '#� i� '#� u� &P� u� &P� i�      >    , �P d� � d� � pl �P pl �P d�      >    , )>� $jD *�� $jD *�� $u� )>� $u� )>� $jD      >    , ��  �X ,�  �X ,�  � ��  � ��  �X      >    , 7� ^� f� ^� f� jL 7� jL 7� ^�      >    , "h�  �� #;�  �� #;�  �8 "h�  �8 "h�  ��      >    , )�� �| *U� �| *U� �4 )�� �4 )�� �|      >    , (�� \ *�� \ *��  (��  (�� \      >    , � &'� �� &'� �� &3L � &3L � &'�      >    , �� 	� �l 	� �l X �� X �� 	�      >    , ې |� 
L |� 
L �D ې �D ې |�      >    , �� !$` Ô !$` Ô !0 �� !0 �� !$`      >    , �P "�4 � "�4 � "�� �P "�� �P "�4      >    , �p #�� �d #�� �d $� �p $� �p #��      >    , r�   T   T � r� � r�        >    , *� � *6� � *6� �� *� �� *� �      >    , !�P 	�� &�( 	�� &�( 
h !�P 
h !�P 	��      >    , '14 � '�� � '�� �� '14 �� '14 �      >    , $�4 |� &  |� &  �D $�4 �D $�4 |�      >    , � ʬ ( ʬ ( �d � �d � ʬ      >    , '�0 	�P )[� 	�P )[� 	� '�0 	� '�0 	�P      >    , ,e< !�L -�P !�L -�P !� ,e< !� ,e< !�L      >    , � ', 	�` ', 	�` 2� � 2� � ',      >    , "�x $C4 "�X $C4 "�X $N� "�x $N� "�x $C4      >    , 
�� %�\   %�\   %� 
�� %� 
�� %�\      >    , } 4 �� 4 �� ?� } ?� } 4      >    , �( � .L � .L �� �( �� �( �      >    , �� 4 Ml 4 Ml ?� �� ?� �� 4      >    , *�� ?t +p ?t +p K, *�� K, *�� ?t      >    , � &'� 2X &'� 2X &3L � &3L � &'�      >    , b� e� �x e� �x q� b� q� b� e�      >    , (�� �� )�L �� )�L �� (�� �� (�� ��      >    , (� !�L )�L !�L )�L !� (� !� (� !�L      >    , #l "� (�� "� (�� "$< #l "$< #l "�      >    , �� �� 	+� �� 	+� �| �� �| �� ��      >    , X $ �H $ �H "� X "� X $      >    , �� =� Z� =� Z� I� �� I� �� =�      >    , � �T �@ �T �@ � � � � �T      >    ,  �� ,� $A@ ,� $A@ 8�  �� 8�  �� ,�      >    , �� e� �� e� �� qh �� qh �� e�      >    , �X !�L vL !�L vL !� �X !� �X !�L      >    , H #�� � #�� � #� H #� H #��      >    , � #�� 0h #�� 0h #ݤ � #ݤ � #��      >    , +�� � -�d � -�d �� +�� �� +�� �      >    , �� �T �� �T �� � �� � �� �T      >    , x %�\ � %�\ � %� x %� x %�\      >    , '� >4 (V, >4 (V, I� '� I� '� >4      >    , �� ( 	�� ( 	�� � �� � �� (      >    , �D �| Y� �| Y� �4 �D �4 �D �|      >    , �� i� 	V� i� 	V� u� �� u� �� i�      >    , J0 #�� cp #�� cp #�| J0 #�| J0 #��      >    , $y� [ 'yx [ 'yx f� $y� f� $y� [      >    , !� �L 8� �L 8� � !� � !� �L      >    , ( < |� (�� |� (�� �D ( < �D ( < |�      >    , #�D =� $� =� $� I� #�D I� #�D =�      >    , ֬ �8 �T �8 �T � ֬ � ֬ �8      >    , )� ( )�� ( )�� � )� � )� (      >    , �4 !�\ � !�\ � " �4 " �4 !�\      >    , �� � �� � �� �� �� �� �� �      >    , -�� �T .�h �T .�h � -�� � -�� �T      >    , %< �8 %�� �8 %�� �� %< �� %< �8      >    , ( !�\ V� !�\ V� " ( " ( !�\      >    , -� �\ .�| �\ .�| � -� � -� �\      >    , Ј �� "($ �� "($ �t Ј �t Ј ��      >    , )�H Đ *DP Đ *DP �H )�H �H )�H Đ      >    , !,0 Wx %ϰ Wx %ϰ c0 !,0 c0 !,0 Wx      >    , !*< D� "� D� "� PX !*< PX !*< D�      >    , �� � #H � #H +� �� +� �� �      >    , L� �\ �T �\ �T � L� � L� �\      >    , �� �P X �P X � �� � �� �P      >    , (<� :l )sT :l )sT F$ (<� F$ (<� :l      >    , �   �   � � � � �        >    , ɐ a| �� a| �� m4 ɐ m4 ɐ a|      >    , .P &l "t &l "t &$ .P &$ .P &l      >    , �( d� !� d� !� p� �( p� �( d�      >    ,  d� �� d� �� p�  p�  d�      >    , 'm� a� '�( a� '�( m� 'm� m� 'm� a�      >    , � $��  �, $��  �, $�L � $�L � $��      >    , 	 � �8 
f �8 
f � 	 � � 	 � �8      >    , (>�   )p   )p � (>� � (>�        >    , %�d %�\ &9( %�\ &9( %� %�d %� %�d %�\      >    , )JP $ )�` $ )�` "� )JP "� )JP $      >    , p( %�d �H %�d �H %� p( %� p( %�d      >    , #� [ $�� [ $�� f� #� f� #� [      >    , �p W0 �H W0 �H b� �p b� �p W0      >    , H� �4 0@ �4 0@ �� H� �� H� �4      >    , 	�D �$ ;  �$ ;  �� 	�D �� 	�D �$      >    , �� =� � =� � I� �� I� �� =�      >    , 	�| � 
 � 
 &| 	�| &| 	�| �      >    , o� 	�P �` 	�P �` 	� o� 	� o� 	�P      >    ,  >4 *� >4 *� I�  I�  >4      >    , O� $"  ~� $"  ~� $-� O� $-� O� $"       >    , �4 %�L � %�L � %� �4 %� �4 %�L      >    , �\ /� ]L /� ]L ;� �\ ;� �\ /�      >    , �4 #�� �D #�� �D #� �4 #� �4 #��      >    , (| �4 (�� �4 (�� �� (| �� (| �4      >    , &�p �� 'q� �� 'q� �D &�p �D &�p ��      >    , ~�    8    8 � ~� � ~�        >    ,  a $פ  �l $פ  �l $�\  a $�\  a $פ      >    , Qt #� �| #� �| /D Qt /D Qt #�      >    , 9 O �� O �� Z� 9 Z� 9 O      >    , �(  �X ��  �X ��  � �(  � �(  �X      >    , � � �@ � �@ h � h � �      >    , %�� �h &` �h &` �  %�� �  %�� �h      >    , �( � � � � �� �( �� �( �      >    , � � Z� � Z� �� � �� � �      >    , �| ;l �� ;l �� G$ �| G$ �| ;l      >    , 4� 7� c� 7� c� C< 4� C< 4� 7�      >    , � �� �@ �� �@ �� � �� � ��      >    , �< � � � � �� �< �� �< �      >    , �� [ �d [ �d f� �� f� �� [      >    , �h %�L ;  %�L ;  %� �h %� �h %�L      >    , zT "� +� "� +� "�� zT "�� zT "�      >    , !7� �� !f� �� !f� �� !7� �� !7� ��      >    , !;� d� "�� d� "�� pl !;� pl !;� d�      >    , v� ', �P ', �P 2� v� 2� v� ',      >    , m� 84 �� 84 �� C� m� C� m� 84      >    , \ d� P d� P p� \ p� \ d�      >    , !�D >4 "�� >4 "�� I� !�D I� !�D >4      >    , B� � � � � �� B� �� B� �      >    , �X !�L �  !�L �  !� �X !� �X !�L      >    , *�� !�L +H !�L +H !� *�� !� *�� !�L      >    , �d !�\ �D !�\ �D " �d " �d !�\      >    , +� �� ,�, �� ,�, �| +� �| +� ��      >    , P � F  � F  �� P �� P �      >    , %0 ʬ %F� ʬ %F� �d %0 �d %0 ʬ      >    , )D �� 0� �� 0� �D )D �D )D ��      >    , $�h   %A   %A � $�h � $�h        >    , U� %�$ O� %�$ O� %�� U� %�� U� %�$      >    , $I ȼ $�� ȼ $�� �t $I �t $I ȼ      >    , �d :l $D :l $D F$ �d F$ �d :l      >    , � �� �� �� �� �| � �| � ��      >    , 'i� #ߘ (�4 #ߘ (�4 #�P 'i� #�P 'i� #ߘ      >    , �0 &l �8 &l �8 &$ �0 &$ �0 &l      >    , W� 	?0 A� 	?0 A� 	J� W� 	J� W� 	?0      >    , � �  �   8 �  8 � �      >    , |(  � 	��  � 	��  � |(  � |(  �      >    , }� � �� � ��  8 }�  8 }� �      >    , �( ��  � ��  � �� �( �� �( ��      >    , �l !$` X� !$` X� !0 �l !0 �l !$`      >    , &� �� ,o  �� ,o  �\ &� �\ &� ��      >    , � |� !l� |� !l� �D � �D � |�      >    , y| \ � \ �  y|  y| \      >    , -� �� .� �� .� � -� � -� ��      >    , f  �� �(  �� �(  �8 f  �8 f  ��      >    ,  0< �� #�� �� #�� ̨  0< ̨  0< ��      >    , %E %�L (� %�L (� %� %E %� %E %�L      >    , v� �4 �$ �4 �$ �� v� �� v� �4      >    , O< O� �� O� �� [� O< [� O< O�      >    , g� JT ,� JT ,� V g� V g� JT      >    , &�( �� '
$ �� '
$ �h &�( �h &�( ��      >    , M�  d ��  d ��  M�  M�  d      >    ,  h x �8 x �8 '0  h '0  h x      >    , �< 
ɸ � 
ɸ � 
�p �< 
�p �< 
ɸ      >    , �X �| 1� �| 1� �4 �X �4 �X �|      >    , 4� [ 6� [ 6� f� 4� f� 4� [      >    , �  ;� R� ;� R� GH �  GH �  ;�      >    , '� i� )� i� )� u� '� u� '� i�      >    , &ό �T 1� �T 1� � &ό � &ό �T      >    , �  d� �  d� �  p� �  p� �  d�      >    , x �8 �@ �8 �@ � x � x �8      >    , $�h  � %�   � %�   �H $�h  �H $�h  �      >    , J !�< � !�< � !�� J !�� J !�<      >    , *|  � *��  � *��  �H *|  �H *|  �      >    , '�� d� (g� d� (g� p� '�� p� '�� d�      >    , x� ~@ �h ~@ �h �� x� �� x� ~@      >    , ]P !�D � !�D � "� ]P "� ]P !�D      >    , &�0 � &�h � &�h �� &�0 �� &�0 �      >    , � �D (� �D (� �� � �� � �D      >    , 5� !�\ /� !�\ /� " 5� " 5� !�\      >    , "W 4 #�@ 4 #�@ ?� "W ?� "W 4      >    , �$ 	X �� 	X ��  �$  �$ 	X      >    , "1� �� $� �� $� �| "1� �| "1� ��      >    , '� !� )�� !� )�� !�� '� !�� '� !�      >    , $�< � &� � &� �� $�< �� $�< �      >    ,  
�h � 
�h � 
�   
�   
�h      >    , 
5H � � � � �X 
5H �X 
5H �      >    , w� �| �� �| �� �4 w� �4 w� �|      >    , ] � � � � �� ] �� ] �      >    ,  � %�$ �8 %�$ �8 %��  � %��  � %�$      >    , 	� �� �� �� �� �� 	� �� 	� ��      >    , "�� #l #x #l #x #"$ "�� #"$ "�� #l      >    , O� 	f@ ( 	f@ ( 	q� O� 	q� O� 	f@      >    , �< %�L C� %�L C� %� �< %� �< %�L      >    , " 
�h �@ 
�h �@ 
�  " 
�  " 
�h      >    , r< � � � � �� r< �� r< �      >    ,  r� � r� � ~d  ~d  r�      >    , !`� 4 !�� 4 !�� ?� !`� ?� !`� 4      >    , � �� W, �� W, �T � �T � ��      >    , � "� �� "� �� "�� � "�� � "�      >    , �0 [ �h [ �h f� �0 f� �0 [      >    , `� "�D `` "�D `` "�� `� "�� `� "�D      >    , $�T �� ._ �� ._ �\ $�T �\ $�T ��      >    , ,��  � -]H  � -]H  � ,��  � ,��  �      >    , �� |� �� |� �� �D �� �D �� |�      >    , �� !�� �h !�� �h !�| �� !�| �� !��      >    ,  � &l � &l � &$  � &$  � &l      >    , �` � @ � @ �� �` �� �` �      >    , �  %�$ �� %�$ �� %�� �  %�� �  %�$      >    , ` � �� � �� �� ` �� ` �      >    , *�� � +>P � +>P �@ *�� �@ *�� �      >    , S� $�� �p $�� �p $�L S� $�L S� $��      >    , &�� ( '�� ( '�� � &�� � &�� (      >    , 4L Đ Θ Đ Θ �H 4L �H 4L Đ      3    , �� �� �D �� �D  ��  �� ��      3    , l` K0 x K0 x �� l` �� l` K0      3    , b� 	�8 nT 	�8 nT 
� b� 
� b� 	�8      3    , m� B� y8 B� y8 �P m� �P m� B�      3    , *8� C� *DP C� *DP �H *8� �H *8� C�      3    , ,i$ � ,t� � ,t� 7� ,i$ 7� ,i$ �      3    , !� � -T � -T � !� � !� �      3    ,  �` &� �` &� �d  �d  �`      3    , )�X � )� � )� 7� )�X 7� )�X �      3    , �0 #۰ �� #۰ �� $�< �0 $�< �0 #۰      3    , �t %�� �, %�� �, &Vt �t &Vt �t %��      3    , G� $�� SD $�� SD %�, G� %�, G� $��      3    , p( 
�� {� 
�� {� �� p( �� p( 
��      3    , �� � � � � �� �� �� �� �      3    , *�h t� *�  t� *�  �t *�h �t *�h t�      3    , '�� �| 'Ť �| 'Ť �� '�� �� '�� �|      3    , )� M� )�H M� )�H �� )� �� )� M�      3    , %Z� 	u� %f8 	u� %f8 	�0 %Z� 	�0 %Z� 	u�      3    , %�� K0 %Ә K0 %Ә �� %�� �� %�� K0      3    , $� 	� $l 	� $l 2� $� 2� $� 	�      3    , %� � %�� � %�� 2� %� 2� %� �      3    , �( �, �� �, �� �T �( �T �( �,      3    , -e Z� -p� Z� -p� �� -e �� -e Z�      3    , X$ J c� J c� ڔ X$ ڔ X$ J      3    , wh �� �  �� �  �� wh �� wh ��      3    , )	� %#� )� %#� )� %� )	� %� )	� %#�      3    ,  � �� � �� I�  I�  �      3    , %C C� %N� C� %N� �� %C �� %C C�   	   3    !    �P  0�  �� 0� $�� +  ,VR_RIGHT_VERTICAL_BUS       3    , *N i, *Y� i, *Y� a *N a *N i,      3    , �� �, �T �, �T o� �� o� �� �,      3    , E0  �0 P�  �0 P� 8� E0 8� E0  �0      3    , q�  ' }h  ' }h  ި q�  ި q�  '      3    , j� � v� � v� �0 j� �0 j� �      3    , $;d J $G J $G �� $;d �� $;d J      3    , )�� �� )�� �� )�� 6� )�� 6� )�� ��      3    , '�� �, '� �, '� H� '�� H� '�� �,      3    , PT �4 \ �4 \ 6� PT 6� PT �4      3    , %n �� %y� �� %y�  %n  %n ��      3    , 
�P %�� 
� %�� 
� &Vt 
�P &Vt 
�P %��      3    , �� � Đ � Đ � �� � �� �      3    , B� � N� � N� �4 B� �4 B� �      3    , ,�� ET -| ET -| �� ,�� �� ,�� ET      3    , ֐ � �H � �H �4 ֐ �4 ֐ �      3    , "Z� J "f� J "f�  � "Z�  � "Z� J      3    , '�� `< '�� `< '�� �l '�� �l '�� `<      3    , E� �� Q� �� Q� 6� E� 6� E� ��      3    , ׬ � �d � �d a ׬ a ׬ �      3    , e$ :l p� :l p� �t e$ �t e$ :l      3    , �X 0� � 0� � :L �X :L �X 0�      3    , 4 \ � \ � 6� 4 6� 4 \      3    , � � �� � ��  �  � �      3    , �� !�� Ь !�� Ь " �� " �� !��      3    , r� $"  ~� $"  ~� %�, r� %�, r� $"       3    , �X %�L � %�L � %�t �X %�t �X %�L      3    , Td �� ` �� ` !t Td !t Td ��      3    ,  �H �  �  �  �  =�  �H =�  �H �      3    , (-( �@ (8� �@ (8� 	bX (-( 	bX (-( �@      3    , 0 �, &� �, &� �4 0 �4 0 �,      3    , � �D H �D H �l � �l � �D      3    ,  6 ��  A� ��  A� Y�  6 Y�  6 ��      3    , �� �� �x �� �x �l �� �l �� ��      3    , ,x !, 80 !, 80 B< ,x B< ,x !,      3    , �� !�� ߜ !�� ߜ "�� �� "�� �� !��      3    , �� �T �d �T �d �4 �� �4 �� �T      3    , ?� �� Kt �� Kt � ?� � ?� ��      3    , �� � �t � �t �� �� �� �� �      3    , K �, V� �, V� N� K N� K �,      3    , )8� � )Dt � )Dt <d )8� <d )8� �      3    , #{� �� #�� �� #�� JX #{� JX #{� ��      3    , �  �� �d  �� �d  ި �  ި �  ��      3    , ��  �� �  �� �  ި ��  ި ��  ��      3    , �l  �T �$  �T �$ �� �l �� �l  �T      3    , y4 i� �� i� �� !� y4 !� y4 i�      3    , r< d� }� d� }� �� r< �� r< d�      3    , -�, �� -�� �� -�� a -�, a -�, ��      3    , ,$� �� ,0� �� ,0� a ,$� a ,$� ��      3    , �� �, �t �, �t  ��  �� �,      3    , �� 	� � 	� � 2� �� 2� �� 	�      3    , $u� C� $�� C� $�� f� $u� f� $u� C�      3    , '�p a� '�( a� '�( � '�p � '�p a�      3    ,  �� ��  �l ��  �l �,  �� �,  �� ��      3    , �� J �� J �� �� �� �� �� J      3    , �P %` � %` � �P �P �P �P %`      3    , �� ^� X ^� X �� �� �� �� ^�      3    , 0�  �� <d  �� <d  ި 0�  ި 0�  ��      3    , #K( h� #V� h� #V� K, #K( K, #K( h�      3    , B �� M� �� M� 6� B 6� B ��      3    , $5�  �0 $A@  �0 $A@ 8� $5� 8� $5�  �0      3    , 
� 28 
� 28 
� 0  
� 0  
� 28      3    , � ~@ �� ~@ �� 7� � 7� � ~@      3    , �� C� � C� � f� �� f� �� C�      3    , %�� 	u� &x 	u� &x 	�0 %�� 	�0 %�� 	u�      3    , )�X �� )� �� )� a )�X a )�X ��      3    , �� |� �� |� �� �� �� �� �� |�      3    , ɔ �� �L �� �L c0 ɔ c0 ɔ ��      3    , �p Ҥ �( Ҥ �( a �p a �p Ҥ      3    , ��  �0 �`  �0 �` �� �� �� ��  �0      3    , �� #� �| #� �| � �� � �� #�      3    , !�$ � !�� � !�� 5� !�$ 5� !�$ �      3    , *ޜ #� *�T #� *�T �4 *ޜ �4 *ޜ #�      3    , '� i� '�H i� '�H � '� � '� i�      3    , '^  �� 'i� �� 'i� 6� '^  6� '^  ��      3    , %�� Ll %�� Ll %�� �� %�� �� %�� Ll      3    , ,| JT ,4 JT ,4 6� ,| 6� ,| JT      3    , �P "� � "� � #�� �P #�� �P "�      3    , �t !�� �, !�� �, "$< �t "$< �t !��      3    , p ]� ( ]� ( �l p �l p ]�      3    , (| t� (+4 t� (+4 �� (| �� (| t�      3    , f� 	u� rd 	u� rd 	� f� 	� f� 	u�      3    , )Y� �0 )e� �0 )e� C� )Y� C� )Y� �0      3    , . t� .� t� .� �� . �� . t�      3    , ,G� _D ,S� _D ,S� a ,G� a ,G� _D      3    , �� K0 ؤ K0 ؤ ٠ �� ٠ �� K0      3    , $�  �� 0�  �� 0�  ި $�  ި $�  ��      3    , �l !$` �$ !$` �$ " �l " �l !$`      3    , +�t G� +�, G� +�, p� +�t p� +�t G�      3    , �� `< �� `< �� �l �� �l �� `<      3    , �< � �� � �� �0 �< �0 �< �      3    , 0 � � � � �0 0 �0 0 �      3    , H� � T@ � T@ �� H� �� H� �      3    , �� J �� J �� g4 �� g4 �� J      3    , X "�\  "�\  #�( X #�( X "�\      3    , 	�d � 	� � 	� 0  	�d 0  	�d �      3    , �� � ݈ � ݈ 0  �� 0  �� �      3    , 	-� �� 	9T �� 	9T � 	-� � 	-� ��      3    , � "?� +\ "?� +\ #�� � #�� � "?�      3    , ?P �� K �� K �� ?P �� ?P ��      3    , � �4 L �4 L 6� � 6� � �4      3    , �t �d �, �d �, �4 �t �4 �t �d      3    , �� � � � � �� �� �� �� �      3    , �( C� 
� C� 
� �� �( �� �( C�      3    , x` �� � �� � �� x` �� x` ��      3    , &�P M� &� M� &� p� &�P p� &�P M�      3    , &�l �T &�$ �T &�$ :L &�l :L &�l �T      3    , %n �T %y� �T %y� :L %n :L %n �T      3    , #�4 � #�� � #�� B@ #�4 B@ #�4 �      3    , #� 6� #�� 6� #�� :L #� :L #� 6�      3    , L$ �� W� �� W� 6� L$ 6� L$ ��      3    , * 	� 5� 	� 5� �� * �� * 	�      3    , �� !�� �\ !�� �\ "�� �� "�� �� !��      3    , 0 �� ;� �� ;� 	bX 0 	bX 0 ��      3    , &l �X &$ �X &$ �P &l �P &l �X      3    , L$ J W� J W� !�� L$ !�� L$ J      3    , � !�� "P !�� "P " � " � !��      3    , �� �d �` �d �` �� �� �� �� �d      3    , 
�t �d 
, �d 
, �� 
�t �� 
�t �d      3    , Gl C� S$ C� S$ � Gl � Gl C�      3    , r� � ~� � ~� 7� r� 7� r� �      3    , 1< �D <� �D <� �� 1< �� 1< �D      3    , $� �, 0� �, 0� �4 $� �4 $� �,      3    , .� �D :� �D :� �l .� �l .� �D      3    , D0 �D O� �D O� �l D0 �l D0 �D      3    , "M@ �� "X� �� "X� '0 "M@ '0 "M@ ��      3    , �� � �� � �� �P �� �P �� �      3    , %)� J %5d J %5d m4 %)� m4 %)� J      3    , ,� !�< 88 !�< 88 !�d ,� !�d ,� !�<      3    , s4 	�P ~� 	�P ~� �� s4 �� s4 	�P      3    , l !�< #$ !�< #$ !�d l !�d l !�<      3    , ')d =� '5 =� '5 a ')d a ')d =�      3    , "tP � "� � "� �� "tP �� "tP �      3    , �4 �< �� �< �� 3, �4 3, �4 �<      3    , 
 � �, 
D �, 
D � 
 � � 
 � �,      3    , 	#� �� 	/� �� 	/� �� 	#� �� 	#� ��      3    , %� �P %H �P %H � %� � %� �P      3    , 4� � @� � @� �0 4� �0 4� �      3    , %� �� %�� �� %�� �� %� �� %� ��      3    , �� �  �\ �  �\ _� �� _� �� �       3    , �� M� �� M� �� �$ �� �$ �� M�      3    , *>t K0 *J, K0 *J, }� *>t }� *>t K0      3    , �| �� �4 �� �4 !�d �| !�d �| ��      3    , Hd $jD T $jD T %�t Hd %�t Hd $jD      3    ,  	, �<  � �<  � !l�  	, !l�  	, �<      3    , �� �< �t �< �t $�< �� $�< �� �<      3    , �� #� а #� а � �� � �� #�      3    , � _  �� _  �� � � � � _       3    , (� � ()@ � ()@ 7� (� 7� (� �      3    , &�< � &�� � &�� �� &�< �� &�< �      3    , %�� � %�H � %�H �� %�� �� %�� �      3    , $�� � %x � %x W� $�� W� $�� �      3    , �  C� � C� � �  �  �  �  C�      3    , �p  �� �(  �� �(  ި �p  ި �p  ��      3    , -�X �� -� �� -� � -�X � -�X ��      3    , �� !� �� !� �� !�d �� !�d �� !�      3    , 80 �� C� �� C� �� 80 �� 80 ��      3    , �� d� Ǡ d� Ǡ �� �� �� �� d�      3    , !�  K0 !�� K0 !�� 
o� !�  
o� !�  K0      3    ,  �  C�  �� C�  �� �X  �  �X  �  C�      3    , -p �� -( �� -( �� -p �� -p ��      3    , ., �� 9� �� 9� VT ., VT ., ��      3    , &�X � &� � &� �p &�X �p &�X �      3    , �� C� �d C� �d �, �� �, �� C�      3    , � �, �` �, �` �4 � �4 � �,      3    , `� Ӝ l` Ӝ l` �� `� �� `� Ӝ      3    , $X� �D $dh �D $dh �l $X� �l $X� �D      3    ,  C� c�  O| c�  O| ��  C� ��  C� c�      3    , �t !� �, !� �, !�d �t !�d �t !�      3    , -A� �� -M� �� -M�  -A�  -A� ��      3    , =� 1 I� 1 I� �P =� �P =� 1      3    , �� 
�h �@ 
�h �@ �� �� �� �� 
�h      3    , � �� | �� | �� � �� � ��      3    , �X �� � �� � �T �X �T �X ��      3    , �l M� �$ M� �$ �t �l �t �l M�      3    , �D � �� � �� 7� �D 7� �D �      3    , !  	u� !� 	u� !� 
L� !  
L� !  	u�      3    ,  � i� ,� i� ,� �  � �  � i�      3    , b� 	u� nT 	u� nT 	� b� 	� b� 	u�      3    , N< x� Y� x� Y� �� N< �� N< x�      3    , x� � �� � �� �\ x� �\ x� �      3    , #� � #< � #< X$ #� X$ #� �      3    , �, J �� J �� �� �, �� �, J      3    , 	�� #�t 	�l #�t 	�l %�� 	�� %�� 	�� #�t      3    , �4 �� �� �� �� �| �4 �| �4 ��      3    , -$� � -0\ � -0\ 	bX -$� 	bX -$� �      3    , &� M� 2� M� 2� �4 &� �4 &� M�      3    , �< �| �� �| �� a �< a �< �|      3    ,  #=|  � #=|  � #��  #��  #=|      3    , !, � ,� � ,� V !, V !, �      3    , *s0 !0 *~� !0 *~� a *s0 a *s0 !0      3    , ip � u( � u( <d ip <d ip �      3    , �  �0 ��  �0 �� 8� � 8� �  �0      3    ,  �  �0  ��  �0  �� 8�  � 8�  �  �0      3    , .p �L :( �L :( :L .p :L .p �L      3    ,  "�� � "�� � #��  #��  "��      3    , %�( �� %�� �� %�� !�@ %�( !�@ %�( ��      3    , (�� �X (� �X (� �P (�� �P (�� �X      3    , )X �d )+ �d )+ �l )X �l )X �d      3    , (� �, (�l �, (�l � (� � (� �,      3    , &�( �, &�� �, &�� � &�( � &�( �,      3    , U| K0 a4 K0 a4 jL U| jL U| K0      3    , � �P �� �P �� � � � � �P      3    , � �� �� �� �� �� � �� � ��      3    , \� t� h� t� h� < \� < \� t�      3    , M$ �� X� �� X� �� M$ �� M$ ��      3    , p( %�D {� %�D {� &$ p( &$ p( %�D      3    , M$ 	?0 X� 	?0 X� 	h4 M$ 	h4 M$ 	?0      3    , � 	?0 &8 	?0 &8 	bX � 	bX � 	?0      3    , tT Đ � Đ � 7� tT 7� tT Đ      3    , L� t� XH t� XH � L� � L� t�      3    , #� #� #H #� #H �L #� �L #� #�      3    , �t  �,  �, a �t a �t       3    , #{� B� #�� B� #�� �� #{� �� #{� B�      3    , + !�� 6� !�� 6� " + " + !��      3    , � !�� � !�� � " � " � !��      3    , �� ~� ߜ ~� ߜ !�d �� !�d �� ~�      3    , xd 	?0 � 	?0 � 	bX xd 	bX xd 	?0      3    , � K0 &8 K0 &8 hX � hX � K0      3    , �T $  � $  � $N� �T $N� �T $       3    , � � l � l F � F � �      3    , � a� < a� < �P � �P � a�      3    , PX F� \ F� \ � PX � PX F�      3    , �  �d �� �d �� �p �  �p �  �d      3    ,  �P �  � �  � �4  �P �4  �P �      3    , O� � [X � [X ,� O� ,� O� �      3    , *�� �� *�x �� *�x a *�� a *�� ��      3    , #�� #�t #�@ #�t #�@ $� #�� $� #�� #�t      3    , !� #�t !�t #�t !�t $� !� $� !� #�t      3    , *�� �d *�H �d *�H K, *�� K, *�� �d      3    , 	�� 	u� 	�� 	u� 	�� 	� 	�� 	� 	�� 	u�      3    , �  	u� �� 	u� �� 	� �  	� �  	u�      3    , �T !� � !� � !�d �T !�d �T !�      3    , � \ �� \ �� D � D � \      3    , 	D J 	� J 	� �T 	D �T 	D J      3    , u( �� �� �� �� a u( a u( ��      3    , 	� M� t M� t �� 	� �� 	� M�      3    ,  �< 	j(  �� 	j(  �� 	�@  �< 	�@  �< 	j(      3    , &+| �D &74 �D &74 �l &+| �l &+| �D      3    , &�  �D &�� �D &�� �l &�  �l &�  �D      3    , �P #�t � #�t � $� �P $� �P #�t      3    , l  Ĭ #$  Ĭ #$ !�0 l !�0 l  Ĭ      3    , *N �$ *Y� �$ *Y� @( *N @( *N �$      3    , #�D =� #�� =� #�� a #�D a #�D =�      3    , R� %�L ^H %�L ^H %�t R� %�t R� %�L      3    ,  d� ?t  p� ?t  p� �T  d� �T  d� ?t      3    , "� Ӝ .l Ӝ .l �l "� �l "� Ӝ      3    , +�4 H +�� H +�� �� +�4 �� +�4 H      3    , �  �T �� �T �� 6� �  6� �  �T      3    , �< H �� H �� :L �< :L �< H      3    , 
A  � 
L� � 
L� � 
A  � 
A  �      3    , U| C� a4 C� a4 �� U| �� U| C�      3    , !;� d� !G� d� !G� �� !;� �� !;� d�      3    , &5@ ET &@� ET &@� nX &5@ nX &5@ ET      3    , �� O� ɐ O� ɐ 0  �� 0  �� O�      3    , 	�D � 	�� � 	�� �� 	�D �� 	�D �      3    , \� � h� � h� �l \� �l \� �      3    , �� �, �\ �, �\ +� �� +� �� �,      3    , � !�� (� !�� (� " � " � !��      3    , �H �d �  �d �  � �H � �H �d      3    , f� K0 r� K0 r� �t f� �t f� K0      3    , �l �� �$ �� �$ %� �l %� �l ��      3    ,   Ll  � Ll  � 6�   6�   Ll      3    , �� "� �� "� �� #�� �� #�� �� "�      3    , k� �� w@ �� w@ �� k� �� k� ��      3    ,  h ��   ��   '0  h '0  h ��      3    , �� x �8 x �8 F �� F �� x      3    , 4 J � J � A� 4 A� 4 J      3    , !A� �4 !Md �4 !Md 6� !A� 6� !A� �4      3    , .4 �� .� �� .� �\ .4 �\ .4 ��      3    , -| D0 -4 D0 -4 ֬ -| ֬ -| D0      3    , b !� m� !� m� !�d b !�d b !�      3    , �P "�4 � "�4 � #�� �P #�� �P "�4      3    , , !�( '� !�( '� "nt , "nt , !�(      3    , .K� �| .WH �| .WH �� .K� �� .K� �|      3    , �� >T �� >T �� �l �� �l �� >T      3    , #� ȼ #�� ȼ #�� a #� a #� ȼ      3    , � � �� � �� 7� � 7� � �      3    , 7� J C� J C� m4 7� m4 7� J      3    ,   !$` � !$` � !�d   !�d   !$`      3    , �,  �� ��  �� ��  ި �,  ި �,  ��      3    , "~ t� "�� t� "�� pl "~ pl "~ t�      3    , �@ $ �� $ �� :L �@ :L �@ $      3    , !j� M� !vh M� !vh p� !j� p� !j� M�      3    , $�  
� $�� 
� $�� � $�  � $�  
�      3    , #+� a\ #7� a\ #7� a #+� a #+� a\      3    , �� � Ԕ � Ԕ �0 �� �0 �� �      3    , � � �� � �� �0 � �0 � �      3    , 
��  �0  h  �0  h X 
�� X 
��  �0      3    , �� �| �� �| �� � �� � �� �|      3    , Fl t� R$ t� R$ G� Fl G� Fl t�      3    , #Ad \ #M \ #M 6� #Ad 6� #Ad \      3    , p� �, |L �, |L d p� d p� �,      3    , �  � �  � � 2� � 2� �  �      3    , 4 � ?� � ?� 2� 4 2� 4 �      3    , �l �, �$ �, �$ �� �l �� �l �,      3    , ,| �� ,4 �� ,4 !�d ,| !�d ,| ��      3    , �� 84 �� 84 �� a �� a �� 84      3    , �� \ �P \ �P 6� �� 6� �� \      3    , !, �� !� �� !� �0 !, �0 !, ��      3    , h ��   ��   �0 h �0 h ��      3    , �  �0 ��  �0 �� �� � �� �  �0      3    , d C�  C�  � d � d C�      3    , �h zX �  zX �  �� �h �� �h zX      3    , 0� K0 <� K0 <� pL 0� pL 0� K0      3    , :� K0 F� K0 F� pL :� pL :� K0      3    , k� ո wD ո wD 	bX k� 	bX k� ո      3    , �L �� � �� � �x �L �x �L ��      3    , �t �� �, �� �, 1 �t 1 �t ��      3    , #t, i� #� i� #� � #t, � #t, i�      3    , !�� i� !� i� !� � !�� � !�� i�      3    , C� � O� � O� 2� C� 2� C� �      3    , > [| I� [| I� �� > �� > [|      3    , �� �| �T �| �T �� �� �� �� �|      3    , &�< C� &�� C� &�� �p &�< �p &�< C�      3    , �| � �4 � �4 oL �| oL �| �      3    ,  f� �  r� �  r� ��  f� ��  f� �      3    , ', 
( 2� 
( 2� �  ', �  ', 
(      3    , "� � "` � "` 6� "� 6� "� �      3    , !�� qh !� qh !� �P !�� �P !�� qh      3    , �� #ټ �t #ټ �t $� �� $� �� #ټ      3    , j� !� v� !� v� !�d j� !�d j� !�      3    , 
P� �� 
\X �� 
\X 
� 
P� 
� 
P� ��      3    , 
s� K0 
� K0 
� �� 
s� �� 
s� K0      3    , "�� � "�� � "�� 7� "�� 7� "�� �      3    , �� J �t J �t ڔ �� ڔ �� J      3    , e� ";� qd ";� qd #�� e� #�� e� ";�      3    , 4� Đ @� Đ @� C` 4� C` 4� Đ      3    , "�� �� "�@ �� "�@  "��  "�� ��      3    , 	H� �< 	T� �< 	T� !0 	H� !0 	H� �<      3    , 	H� 8T 	T� 8T 	T� �� 	H� �� 	H� 8T      3    , Wp � c( � c( �� Wp �� Wp �      3    , _D 
= j� 
= j� � _D � _D 
=      3    , i0 K0 t� K0 t� �� i0 �� i0 K0      3    , �$ $ �� $ �� :L �$ :L �$ $      3    , �� M� �� M� �� �$ �� �$ �� M�      3    , �  � � � � �4 �  �4 �  �      3    , � >4 *d >4 *d j� � j� � >4      3    , 	�| M� 	�4 M� 	�4 &| 	�| &| 	�| M�      3    , Fp � R( � R( �4 Fp �4 Fp �      3    , �� �, �� �, �� �T �� �T �� �,      3    , d� t� pl t� pl �� d� �� d� t�      3    , �< %�L �� %�L �� %�t �< %�t �< %�L      3    , \� %�  hT %�  hT &$ \� &$ \� %�       3    , "�\ r� "� r� "� ;� "�\ ;� "�\ r�      3    , ?P � K � K � ?P � ?P �      3    , %�� �� %�� �� %��  %��  %�� ��      3    , ,2t �< ,>, �< ,>, �� ,2t �� ,2t �<      3    , � �� �P �� �P �� � �� � ��      3    , �� �� �h �� �h �� �� �� �� ��      3    , l  �0 $  �0 $ X l X l  �0      3    , �P  �0 �  �0 � X �P X �P  �0      3    ,  �� ��  �� ��  �� /D  �� /D  �� ��      3    , R  t� ]� t� ]� �� R  �� R  t�      3    , P � ' � ' �� P �� P �      3    , 	h4 � 	s� � 	s� < 	h4 < 	h4 �      3    , 	#� ` 	/� ` 	/� < 	#� < 	#� `      3    , �� �< ̤ �< ̤ !W( �� !W( �� �<      3    , �d "l � "l � #�� �d #�� �d "l      3    , 3� J ?t J ?t �\ 3� �\ 3� J      3    , %�� =� %�� =� %�� � %�� � %�� =�      3    , Y  �  d� �  d� � Y  � Y  �       3    , �� � ܈ � ܈ �4 �� �4 �� �      3    , �, 
`@ �� 
`@ �� � �, � �, 
`@      3    , #� 	u� /H 	u� /H 
k� #� 
k� #� 	u�      3    , �� C� 	� C� 	� �� �� �� �� C�      3    , D �� � �� � ?� D ?� D ��      3    , �X �d � �d � �� �X �� �X �d      3    , �H �d   �d   �� �H �� �H �d      3    , � "� +� "� +� #�� � #�� � "�      3    , #9� !�4 #EL !�4 #EL "�� #9� "�� #9� !�4      3    , �� U| ܬ U| ܬ �� �� �� �� U|      3    , �D M� �� M� �� l� �D l� �D M�      3    , !G� ȼ !S@ ȼ !S@ l� !G� l� !G� ȼ      3    , �� � ۔ � ۔ @L �� @L �� �      3    , �� 4� �8 4� �8 a �� a �� 4�      3    , �, $f\ �� $f\ �� %�t �, %�t �, $f\      3    , 
� #�t 
#� #�t 
#� $+� 
� $+� 
� #�t      3    ,  | M� ,4 M� ,4 �L  | �L  | M�      3    , �� �d � �d � � �� � �� �d      3    , 3� �| ?x �| ?x �� 3� �� 3� �|      3    , � �� �t �� �t �� � �� � ��      3    , "� U| "�\ U| "�\ �� "� �� "� U|      3    , .� �� :H �� :H � .� � .� ��      3    , �, �� �� �� �� � �, � �, ��      3    , $�� �� $�d �� $�d @ $�� @ $�� ��      3    , 
h "� 
s� "� 
s� #�� 
h #�� 
h "�      3    , -�p �d .	( �d .	( �� -�p �� -�p �d      3    , K, t� V� t� V� �� K, �� K, t�      3    , $� t� $�� t� $�� �< $� �< $� t�      3    , 1� 	u� =� 	u� =� 
�H 1� 
�H 1� 	u�      3    , zx 
�� �0 
�� �0 � zx � zx 
��      3    , |$ K0 �� K0 �� C< |$ C< |$ K0      3    , � � l � l � � � � �      3    , _� �L kh �L kh :L _� :L _� �L      3    , �� 	u� �` 	u� �` 	� �� 	� �� 	u�      3    , � 	u� &8 	u� &8 #  � #  � 	u�      3    , .P ?x : ?x : �� .P �� .P ?x      3    , �� C� � C� � f� �� f� �� C�      3    , � %�� 8 %�� 8 &$ � &$ � %��      3    , 	� L 	8 L 	8 �� 	� �� 	� L      3    , 	�@ �d 	�� �d 	�� ( 	�@ ( 	�@ �d      3    , #\� |� #ht |� #ht �� #\� �� #\� |�      3    , $`� |� $l8 |� $l8 �� $`� �� $`� |�      3    , _D 	?0 j� 	?0 j� 	bX _D 	bX _D 	?0      3    , Kt �� W, �� W, a Kt a Kt ��      3    , ֈ  d �@  d �@ �4 ֈ �4 ֈ  d      3    , '� K0 '#� K0 '#� 	� '� 	� '� K0      3    , b� � n| � n| �� b� �� b� �      3    , �H 6� �  6� �  p� �H p� �H 6�      3    , Q � \� � \� B@ Q B@ Q �      3    , �� d� �h d� �h �� �� �� �� d�      3    , oL �d { �d { �� oL �� oL �d      3    , 
�� d� 
�H d� 
�H �� 
�� �� 
�� d�      3    , 
�8 t 
�� t 
�� B< 
�8 B< 
�8 t      3    , �� �@ �� �@ ��  ��  �� �@      3    , }� � �� � �� 7� }� 7� }� �      3    , zT !�� � !�� � #"$ zT #"$ zT !��      3    , �8 84 �� 84 �� �� �8 �� �8 84      3    , �` �� � �� � a �` a �` ��      3    , \� � hT � hT 	bX \� 	bX \� �      3    , x� � �� � �� 0  x� 0  x� �      3    , u, C� �� C� �� �X u, �X u, C�      3    , 2� � >� � >� 7� 2� 7� 2� �      3    , � !�< %� !�< %� !�@ � !�@ � !�<      3    , �� !�� �� !�� �� " �� " �� !��      3    , �| v� �4 v� �4 @( �| @( �| v�      3    , S� d� _h d� _h �� S� �� S� d�      3    , e� �d q� �d q� �4 e� �4 e� �d      3    , �H �, �  �, �  �T �H �T �H �,      3    , �� �, �d �, �d q� �� q� �� �,      3    , �4 ٜ �� ٜ �� �$ �4 �$ �4 ٜ      3    , !� �L !�h �L !�h �� !� �� !� �L      3    , "&0 M� "1� M� "1� � "&0 � "&0 M�      3    , *�( �, *�� �, *�� �� *�( �� *�( �,      3    , m� � y8 � y8 "� m� "� m� �      3    , K0 !�� V� !�� V� " K0 " K0 !��      3    , ( ed 3� ed 3� " ( " ( ed      3    , *4� �� *@h �� *@h �� *4� �� *4� ��      3    , � �d %� �d %� K, � K, � �d      3    , �4 ٜ �� ٜ �� �l �4 �l �4 ٜ      3    ,  0< C�  ;� C�  ;� �H  0< �H  0< C�      3    ,  �D K0  �� K0  �� hX  �D hX  �D K0      3    , � D0 �� D0 �� �\ � �\ � D0      3    , _� 	p k@ 	p k@ #  _� #  _� 	p      3    , �� H �h H �h :L �� :L �� H      3    , �| #l �4 #l �4 #�� �| #�� �| #l      3    , �4 J �� J �� ڔ �4 ڔ �4 J      3    , �� J � J � �l �� �l �� J      3    , 	�0 f< 	�� f< 	�� �l 	�0 �l 	�0 f<      3    , D �d � �d � �� D �� D �d      3    , �� H �x H �x F �� F �� H      3    , t t� ", t� ", $d t $d t t�      3    , \4 � g� � g� �l \4 �l \4 �      3    , :� �l FL �l FL �\ :� �\ :� �l      3    , �� #�t �` #�t �` $� �� $� �� #�t      3    , SH �( _  �( _  �P SH �P SH �(      3    , Gl �( S$ �( S$ �P Gl �P Gl �(      3    , p 	u� ( 	u� ( 	�` p 	�` p 	u�      3    , #Z� C� #f� C� #f� �p #Z� �p #Z� C�      3    , �� "b� �l "b� �l #�� �� #�� �� "b�      3    , "* �� "5� �� "5� ct "* ct "* ��      3    , )[� �< )g� �< )g� �d )[� �d )[� �<      3    , (�� J (� J (� �� (�� �� (�� J      3    , 4P $�l @ $�l @ %�, 4P %�, 4P $�l      3    , �� #�t �\ #�t �\ $�$ �� $�$ �� #�t      3    , _� �� k� �� k� � _� � _� ��      3    , �� �� �� �� �� � �� � �� ��      3    , ݬ #�t �d #�t �d $/� ݬ $/� ݬ #�t      3    , �� �� Ҥ �� Ҥ 6� �� 6� �� ��      3    , �( �d �� �d �� � �( � �( �d      3    , R� K0 ^� K0 ^� �� R� �� R� K0      3    , )H �� 5  �� 5  	h4 )H 	h4 )H ��      3    , !7� �� !C� �� !C� �� !7� �� !7� ��      3    , -�( �, -�� �, -�� �T -�( �T -�( �,      3    , >� 	 J� 	 J� 	bX >� 	bX >� 	      3    , 	�x 	 	�0 	 	�0 	bX 	�x 	bX 	�x 	      3    , ,0� �� ,<8 �� ,<8 u� ,0� u� ,0� ��      3    , �� �� �� �� �� m� �� m� �� ��      3    , *B\ � *N � *N 7� *B\ 7� *B\ �      3    , )�X {� )� {� )� 	n )�X 	n )�X {�      3    , �< ^� �� ^� �� fd �< fd �< ^�      3    , �L 	u� � 	u� � 
H� �L 
H� �L 	u�      3    , P �� ' �� ' �8 P �8 P ��      3    , *�� �� *�� �� *�� �� *�� �� *�� ��      3    , �� i� �h i� �h � �� � �� i�      3    , �� �� �� �� �� ø �� ø �� ��      3    , �� $ � �8 $ � �8 %�t �� %�t �� $ �      3    , G$ �< R� �< R� !0 G$ !0 G$ �<      3    ,  � 
ɸ � 
ɸ � �  � �  � 
ɸ      3    , ې � �H � �H �4 ې �4 ې �      3    , M� �| Y� �| Y� �� M� �� M� �|      3    , -ΐ � -�H � -�H F -ΐ F -ΐ �      3    , �( �( �� �( �� �0 �( �0 �( �(      3    , 
�� t� 
�� t� 
�� �� 
�� �� 
�� t�      3    , ,�� �` ,�� �` ,�� !� ,�� !� ,�� �`      3    , #t, t� #� t� #� �� #t, �� #t, t�      3    , �� �(  � �(  � � �� � �� �(      3    , �@ M� �� M� �� a �@ a �@ M�      3    , �� $ �8 $ �8 :L �� :L �� $      3    , � !�< *� !�< *� !�d � !�d � !�<      3    , �� � �t � �t 2� �� 2� �� �      3    , /� � ;h � ;h 2� /� 2� /� �      3    , �< \� � \� � 	n �< 	n �< \�      3    , %�l �� %�$ �� %�$ �� %�l �� %�l ��      3    , #�� �d #�l �d #�l �| #�� �| #�� �d      3    , �0 !�< �� !�< �� !�d �0 !�d �0 !�<      3    , ې |� �H |� �H �� ې �� ې |�      3    , �� � �H � �H 7� �� 7� �� �      3    , �� �P 	x �P 	x �$ �� �$ �� �P      3    , 
7<  
B�  
B� 2� 
7< 2� 
7<       3    , &ɰ !�� &�h !�� &�h " &ɰ " &ɰ !��      3    , #� !�� #ټ !�� #ټ "j� #� "j� #� !��      3    , �| t� �4 t� �4 �� �| �� �| t�      3    , �� G� �L G� �L a �� a �� G�      3    , $�� Đ $٘ Đ $٘ 7� $�� 7� $�� Đ      3    , ,G� �@ ,S� �@ ,S� 	bX ,G� 	bX ,G� �@      3    , 	T �  �  =� 	T =� 	T �      3    , � C� �� C� �� �p � �p � C�      3    , 2x %�D >0 %�D >0 &3L 2x &3L 2x %�D      3    , ,�� �  -| �  -| @L ,�� @L ,�� �       3    , ,o  4� ,z� 4� ,z� :L ,o  :L ,o  4�      3    , �� �4 �� �4 �� �� �� �� �� �4      3    , B� $ N� $ N� :L B� :L B� $      3    , 
�@ �, 
�� �, 
�� �4 
�@ �4 
�@ �,      3    , �T !�< � !�< � !�d �T !�d �T !�<      3    , �P |� � |� � �� �P �� �P |�      3    , l Z� w� Z� w� 	bX l 	bX l Z�      3    , � C� �@ C� �@ �H � �H � C�      3    , 
1` G� 
= G� 
= ?� 
1` ?� 
1` G�      3    , �p �| �( �| �( �� �p �� �p �|      3    , � 	?0 � 	?0 � 	bX � 	bX � 	?0      3    , �H t� �  t� �  $d �H $d �H t�      3    , !� b� -� b� -� �� !� �� !� b�      3    , J �� U� �� U� �� J �� J ��      3    , �h A� �  A� �  �� �h �� �h A�      3    , #(  d� #3� d� #3� �� #(  �� #(  d�      3    , �� :l �8 :l �8 �� �� �� �� :l      3    , �l �$ �$ �$ �$ �� �l �� �l �$      3    , %�h �� %�  �� %�  �0 %�h �0 %�h ��      3    , |  � &4  � &4 8� | 8� |  �      3    , '� � '�� � '�� �� '� �� '� �      3    , '14 t� '<� t� '<� �� '14 �� '14 t�      3    , �H |� �  |� �  �� �H �� �H |�      3    , !� W� !� W� !� :L !� :L !� W�      3    , P %��  %��  &$ P &$ P %��      3    , �, %�� �� %�� �� &$ �, &$ �, %��      3    , �� �� ƨ �� ƨ ø �� ø �� ��      3    , �l K0 �$ K0 �$   �l   �l K0      3    , �0 \ �� \ �� 	bX �0 	bX �0 \      3    , x� �� �@ �� �@ 	bX x� 	bX x� ��      3    , �� � �l � �l < �� < �� �      3    , � �, � �, � �T � �T � �,      3    , �0 ٜ �� ٜ �� �l �0 �l �0 ٜ      3    , '/@ �� ':� �� ':�  '/@  '/@ ��      3    , �T ,� � ,� � � �T � �T ,�      3    , � ( L ( L 4, � 4, � (      3    , ��  �0 �  �0 � �� �� �� ��  �0      3    , �� �, � �, � �T �� �T �� �,      3    , 
� C� 
�� C� 
�� �  
� �  
� C�      3    , ._ #�t .j� #�t .j� $R� ._ $R� ._ #�t      3    , )mx $G )y0 $G )y0 %�� )mx %�� )mx $G      3    , "� �� "� �� "� �8 "� �8 "� ��      3    , 5h #۰ A  #۰ A  $� 5h $� 5h #۰      3    , �� #�t �� #�t �� $� �� $� �� #�t      3    , !Kp 	?0 !W( 	?0 !W( 	bX !Kp 	bX !Kp 	?0      3    , 	��  �0 	�`  �0 	�` _� 	�� _� 	��  �0      3    , �h �< �  �< �  !�� �h !�� �h �<      3    , .� � :L � :L �4 .� �4 .� �      3    , "5� !�< "A� !�< "A� !�d "5� !�d "5� !�<      3    , !n�  Ĭ !zP  Ĭ !zP !�0 !n� !�0 !n�  Ĭ      3    , (�� � (�� � (�� �0 (�� �0 (�� �      3    ,  _ �  j� �  j� 7�  _ 7�  _ �      3    , &�l 6� &�$ 6� &�$ �H &�l �H &�l 6�      3    , #�� � $� � $� �� #�� �� #�� �      3    , w� �| �� �| �� �� w� �� w� �|      3    , �� �| �� �| �� �$ �� �$ �� �|      3    , )l >T 5$ >T 5$ iL )l iL )l >T      3    , � �, +� �, +� +� � +� � �,      3    , !�< �� !�� �� !�� 	bX !�< 	bX !�< ��      3    , !� C� !� C� !� f� !� f� !� C�      3    , "� C� "�� C� "�� f� "� f� "� C�      3    , #� �, #H �, #H +� #� +� #� �,      3    , +�0 t� +�� t� +�� �� +�0 �� +�0 t�      3    , '�  i� '�� i� '�� �4 '�  �4 '�  i�      3    , uP J � J � �D uP �D uP J      3    , ld J x J x m4 ld m4 ld J      3    , � �< �� �< �� �d � �d � �<      3    , �� \ �P \ �P 6� �� 6� �� \      3    , �� \ �� \ �� 6� �� 6� �� \      3    , g �� r� �� r� ø g ø g ��      3    , �� 	u� �T 	u� �T q� �� q� �� 	u�      3    , r�  �0 ~�  �0 ~� X r� X r�  �0      3    , {P S� � S� � �0 {P �0 {P S�      3    , 
�� \� 
ϔ \� 
ϔ q� 
�� q� 
�� \�      3    , b�  �0 nT  �0 nT X b� X b�  �0      3    , �l �h �$ �h �$ 7� �l 7� �l �h      3    , -�D 	p -�� 	p -�� VX -�D VX -�D 	p      3    , �, w  �� w  �� �0 �, �0 �, w       3    , ]�  �0 iP  �0 iP X ]� X ]�  �0      3    , �4 %�L �� %�L �� %�t �4 %�t �4 %�L      3    , RH �< ^  �< ^   �� RH  �� RH �<      3    , �� $�� �h $�� �h %�t �� %�t �� $��      3    , (!p �d (-( �d (-( �� (!p �� (!p �d      3    , %�� �� %�� �� %�� � %�� � %�� ��      3    , $hP �d $t �d $t � $hP � $hP �d      3    , $�h �� $�  �� $�  �� $�h �� $�h ��      3    , '�( d� '�� d� '�� �� '�( �� '�( d�      3    , 	/� h� 	;H h� 	;H � 	/� � 	/� h�      3    , �L �\  �\  �\ �L �\ �L �\      3    , #nP o� #z o� #z �4 #nP �4 #nP o�      3    , � �� � �� � �p � �p � ��      3    , ] � h� � h� �4 ] �4 ] �      3    , *�� \ *�� \ *�� 6� *�� 6� *�� \      3    , (�� \ (�� \ (�� 6� (�� 6� (�� \      3    , "� �D ""H �D ""H �l "� �l "� �D      3    , .�� �, .�h �, .�h � .�� � .�� �,      3    , #l �� #"$ �� #"$  #l  #l ��      3    , 	\| � 	h4 � 	h4 �4 	\| �4 	\| �      3    , 9P �� E �� E @ 9P @ 9P ��      3    , �h �� �  �� �  @ �h @ �h ��      3    , & [ 1� [ 1� 7� & 7� & [      3    , �� � � � � )  �� )  �� �      3    , +]� Z� +iH Z� +iH �� +]� �� +]� Z�      3    , ϐ �� �H �� �H �X ϐ �X ϐ ��      3    ,  �� d�  � d�  � ��  �� ��  �� d�      3    , )  � )� � )� 0  )  0  )  �      3    , (�� C� (�� C� (�� �  (�� �  (�� C�      3    , �� �� �� �� �� �� �� �� �� ��      3    , "�� Đ "� Đ "� 7� "�� 7� "�� Đ      3    , 4 � � � � �0 4 �0 4 �      3    , �X � � � � 7� �X 7� �X �      3    , �0 M� �� M� �� p� �0 p� �0 M�      3    , r� � ~` � ~` :L r� :L r� �      3    , �� M� �x M� �x I� �� I� �� M�      3    , � � %� � %� �� � �� � �      3    , %0 �< %� �< %� �d %0 �d %0 �<      3    , $0 �< $%� �< $%�  � $0  � $0 �<      3    , �p S� �( S� �( :L �p :L �p S�      3    , x � �� � �� _� x _� x �      3    , $)� ~� $5� ~� $5� l� $)� l� $)� ~�      3    , $�� �T $�� �T $�� �< $�� �< $�� �T      3    , %bP �@ %n �@ %n 	bX %bP 	bX %bP �@      3    , ${� 
ш $�� 
ш $�� � ${� � ${� 
ш      3    , �, [| �� [| �� ~� �, ~� �, [|      3    , �$ %�� �� %�� �� &$ �$ &$ �$ %��      3    , �� s �t s �t �0 �� �0 �� s      3    , 1� 7� =� 7� =� 	bX 1� 	bX 1� 7�      3    , �$ �� �� �� �� hX �$ hX �$ ��      3    , � �d � �d � �| � �| � �d      3    , � � !t � !t �� � �� � �      3    , Yd �� e �� e 	n Yd 	n Yd ��      3    , K0 �� V� �� V� �� K0 �� K0 ��      3    , ¼ � �t � �t �4 ¼ �4 ¼ �      3    , �� [| �x [| �x �� �� �� �� [|      3    , "`� %�� "l� %�� "l� &$ "`� &$ "`� %��      3    ,  a #�t  l� #�t  l� $�\  a $�\  a #�t      3    , �� K0 �@ K0 �@ �t �� �t �� K0      3    , ʰ i� �h i� �h � ʰ � ʰ i�      3    , U� t� a� t� a� �� U� �� U� t�      3    , � =� l =� l a � a � =�      3    , �� "b� �� "b� �� #�� �� #�� �� "b�      3    , !�@ � !�� � !�� 	bX !�@ 	bX !�@ �      3    , !� �h !�� �h !�� �� !� �� !� �h      3    , 	��  � 	��  � 	��  ި 	��  ި 	��  �      3    , �  �� ��  �� ��  ި �  ި �  ��      3    , "l� �� "x8 �� "x8 �� "l� �� "l� ��      3    , 	}� � 	�h � 	�h 7� 	}� 7� 	}� �      3    , ~� � �� � �� 7� ~� 7� ~� �      3    , wh 	u� �  	u� �  	�X wh 	�X wh 	u�      3    , � K0 @ K0 @ �� � �� � K0      3    , -A� �d -M� �d -M� �� -A� �� -A� �d      3    , X�  �0 dH  �0 dH X X� X X�  �0      3    , ƀ #�t �8 #�t �8 $r ƀ $r ƀ #�t      3    , �< $ �� $ �� :L �< :L �< $      3    , �� �< �X �< �X �� �� �� �� �<      3    , +� �4 7� �4 7� 6� +� 6� +� �4      3    , 'VP 8T 'b 8T 'b �� 'VP �� 'VP 8T      3    , &� 8T &�� 8T &�� �� &� �� &� 8T      3    , ��  �x ��  �x �� X �� X ��  �x      3    , _� %�� kd %�� kd &3L _� &3L _� %��      3    , �� |� ڔ |� ڔ �� �� �� �� |�      3    , '� !� '#� !� '#� !�d '� !�d '� !�      3    , }h z� �  z� �  0  }h 0  }h z�      3    , P| � \4 � \4 0  P| 0  P| �      3    , R� � ^H � ^H 0  R� 0  R� �      3    , �� @ Ր @ Ր � �� � �� @      3    , �0 � �� � �� 0  �0 0  �0 �      3    , !� �< ! x �< ! x  �d !�  �d !� �<      3    , +d J + J +  �d +d  �d +d J      3    , �$ K0 �� K0 �� �t �$ �t �$ K0      3    , Ƥ � �\ � �\ g4 Ƥ g4 Ƥ �      3    , #l !�� #"$ !�� #"$ "$< #l "$< #l !��      3    , !�� b� !� b� !� hX !�� hX !�� b�      3    , " K0 "� K0 "� hX " hX " K0      3    , �� *h �t *h �t 0  �� 0  �� *h      3    , ��  �0 ��  �0 �� ~� �� ~� ��  �0      3    , $�| \ $�4 \ $�4 6� $�| 6� $�| \      3    , %�@ \ %�� \ %�� 6� %�@ 6� %�@ \      3    , *�� C� *�H C� *�H �@ *�� �@ *�� C�      3    , {, #�t �� #�t �� $R� {, $R� {, #�t      3    , �@ K0 �� K0 �� fd �@ fd �@ K0      3    , e� �� q@ �� q@ 6  e� 6  e� ��      3    , 4 	u� � 	u� � �� 4 �� 4 	u�      3    , �  �0 ��  �0 �� �� � �� �  �0      3    , �$ !=� �� !=� �� !�d �$ !�d �$ !=�      3    , d J  J  !I| d !I| d J      3    , )0� >� )<� >� )<� �P )0� �P )0� >�      3    , $�� 	 %� 	 %� 	bX $�� 	bX $�� 	      3    , 'VP 	 'b 	 'b 	bX 'VP 	bX 'VP 	      3    , ~� �d �� �d �� �� ~� �� ~� �d      3    , 1�  �0 =�  �0 =� X 1� X 1�  �0      3    , � �� �� �� �� JX � JX � ��      3    ,  (l �d  4$ �d  4$ �  (l �  (l �d      3    , -|� 	u� -�@ 	u� -�@ Rp -|� Rp -|� 	u�      3    , #�� Ӝ #�d Ӝ #�d �l #�� �l #�� Ӝ      3    , 	� t� � t� � �� 	� �� 	� t�      3    , H �� #  �� #  @ H @ H ��      3    , "� K0 .t K0 .t �� "� �� "� K0      3    , -�  �� 9t  �� 9t  ި -�  ި -�  ��      3    , ��  �� �h  �� �h  ި ��  ި ��  ��      3    , &�P #�� &� #�� &� #�� &�P #�� &�P #��      3    , & #�� &� #�� &� #�� & #�� & #��      3    , .� Ӝ :� Ӝ :� �8 .� �8 .� Ӝ      3    , +u  �� +�� �� +�� =� +u  =� +u  ��      3    , (/  �� (:�  �� (:�  ި (/  ި (/  ��      3    , - � -� � -� 7� - 7� - �      3    , +�� ?x +ڐ ?x +ڐ nX +�� nX +�� ?x      3    , �< i, �� i, �� a �< a �< i,      3    , )� �$ 5h �$ 5h :L )� :L )� �$      3    , C� M� O� M� O� p� C� p� C� M�      3    , ��  �� �P  �� �P  ި ��  ި ��  ��      3    , r� �< ~< �< ~< !� r� !� r� �<      3    , ]� _D iP _D iP ?� ]� ?� ]� _D      3    , ~� � �� � �� �� ~� �� ~� �      3    , T K0  K0  �t T �t T K0      3    , a� ^� m8 ^� m8 �t a� �t a� ^�      3    , b #�t m� #�t m� $� b $� b #�t   	   3    !    �  � Q � T�      3    , D � � � � L( D L( D �      3    , < |� $� |� $� �� < �� < |�      3    ,  �p   �(   �( 0   �p 0   �p       3    , 	� S� � S� � :L 	� :L 	� S�      3    , � 	u� �8 	u� �8 	� � 	� � 	u�      3    , �� 	u� �| 	u� �| 	� �� 	� �� 	u�      3    , !,0 Wx !7� Wx !7� C` !,0 C` !,0 Wx      3    , !*< K0 !5� K0 !5� PX !*< PX !*< K0      3    , ( < h (� h (� 	bX ( < 	bX ( < h      3    , (ŀ K0 (�8 K0 (�8   (ŀ   (ŀ K0      3    , (, >X 3� >X 3� :L (, :L (, >X      3    , [< >X f� >X f� :L [< :L [< >X      3    , 
\ � 
 � 
 a 
\ a 
\ �      3    , $� t� 0@ t� 0@ �� $� �� $� t�      3    , ߠ �� �X �� �X B� ߠ B� ߠ ��      3    , q� �  }@ �  }@ �P q� �P q� �       3    , |� �D �L �D �L �l |� �l |� �D      3    , ֬ #�t �d #�t �d $� ֬ $� ֬ #�t      3    , g� %�L s� %�L s� %�t g� %�t g� %�L      3    , �� ~� �X ~� �X �� �� �� �� ~�      3    , �p !�< 
( !�< 
( !�d �p !�d �p !�<      3    , )�| F� )�4 F� )�4 �� )�| �� )�| F�      3    , %H� �� %T� �� %T� �� %H� �� %H� ��      3    , (8� !�� (D� !�� (D� " (8� " (8� !��      3    , &�� !�< &͘ !�< &͘ !�d &�� !�d &�� !�<      3    , %< �  %� �  %� �� %< �� %< �       3    , &�� �  &�� �  &�� � &�� � &�� �       3    , � �� � �� � �0 � �0 � ��      3    , � K0 �H K0 �H fd � fd � K0      3    , �� =� � =� � a �� a �� =�      3    , N� =� Z� =� Z� a N� a N� =�      3    , *�p �� *�( �� *�( : *�p : *�p ��      3    , 'e� �� 'q� �� 'q� ø 'e� ø 'e� ��      3    , 
�< �| 
�� �| 
�� �� 
�< �� 
�< �|      3    , C� �� O� �� O�  8 C�  8 C� ��      3    , m8 
d( x� 
d( x� � m8 � m8 
d(      3    , �� hT �d hT �d �� �� �� �� hT      3    , [� �, g\ �, g\ q� [� q� [� �,      3    , ct hT o, hT o, �� ct �� ct hT      3    , � C� �� C� �� f� � f� � C�      3    , 
 �P � �P � 7� 
 7� 
 �P      3    , $�p a� $�( a� $�( �P $�p �P $�p a�      3    , %h, �d %s� �d %s� �� %h, �� %h, �d      3    , #�� �d #� �d #� �� #�� �� #�� �d      3    , -�4 �� -�� �� -�� �� -�4 �� -�4 ��      3    , -� �� -(� �� -(� F$ -� F$ -� ��      3    , �4 !�� �� !�� �� " �4 " �4 !��      3    , '�� $ '�� $ '�� :L '�� :L '�� $      3    , $t 	�P $� 	�P $� 
�0 $t 
�0 $t 	�P   	   3    !    �  (<� � (<� �      3    , �, �T �� �T �� �� �, �� �, �T      3    , �� $ �� $ �� :L �� :L �� $      3    ,  f�  �X  r�  �X  r�  ި  f�  ި  f�  �X      3    , � C�  X C�  X �H � �H � C�      3    , �< \ �� \ �� B< �< B< �< \      3    , *4� � *@h � *@h )  *4� )  *4� �      3    , *�� � *ܨ � *ܨ )  *�� )  *�� �      3    , � �� �� �� ��  �  � ��      3    , ', �� 2� �� 2�  ',  ', ��      3    , )� $ )�` $ )�` :L )� :L )� $      3    , +K� t� +W� t� +W� �� +K� �� +K� t�      3    , �@ �< �� �< �� !W( �@ !W( �@ �<      3    , �| �l �4 �l �4 a �| a �| �l      3    , *| \� *4 \� *4 
� *| 
� *| \�      3    , %�� 	u� %׀ 	u� %׀ 
�@ %�� 
�@ %�� 	u�      3    , �� �� ֈ �� ֈ �, �� �, �� ��      3    , �� !�< ` !�< ` !�d �� !�d �� !�<      3    , W �, b� �, b� | W | W �,      3    , x� C� �@ C� �@ �� x� �� x� C�      3    , ��  �� ˈ  �� ˈ  ި ��  ި ��  ��      3    , �p  �� �(  �� �(  ި �p  ި �p  ��      3    , �0  �� �  �� �  ި �0  ި �0  ��      3    , (0 !�� (�� !�� (�� "$< (0 "$< (0 !��      3    , (�� !�� (ŀ !�� (ŀ "j� (�� "j� (�� !��      3    , *p b� *!( b� *!( hX *p hX *p b�      3    , )�� K0 )�8 K0 )�8 hX )�� hX )�� K0      3    , (c� �d (o� �d (o� � (c� � (c� �d      3    , $E( �d $P� �d $P� � $E( � $E( �d      3    , .�  �0 :�  �0 :� X .� X .�  �0      3    , R � ]� � ]� �0 R �0 R �      3    , �, C� �� C� �� C` �, C` �, C�      3    , q� � }h � }h @ q� @ q� �      3    , dH 	u� p  	u� p  
h dH 
h dH 	u�      3    , < $f\ � $f\ � %�t < %�t < $f\      3    , ,� C� 8� C� 8� �  ,� �  ,� C�      3    , �� � � � � 0  �� 0  �� �      3    , � 	j( � 	j( � 	� � 	� � 	j(      3    , �� �  �P �  �P �P �� �P �� �       3    , �4 �d �� �d �� �4 �4 �4 �4 �d      3    , z� �| �� �| �� �� z� �� z� �|      3    , $�h �� $�  �� $�  �� $�h �� $�h ��      3    , & � F� &< F� &< � & � � & � F�      3    , { 	u� �� 	u� �� 
� { 
� { 	u�      3    , ,�� �D ,�� �D ,�� �l ,�� �l ,�� �D      3    ,  Ĭ ��  �d ��  �d :L  Ĭ :L  Ĭ ��      3    , |� �� �h �� �h :L |� :L |� ��      3    , m� t� yX t� yX �� m� �� m� t�      3    , k� t� w@ t� w@ �� k� �� k� t�      3    , +q #�t +|� #�t +|� %�, +q %�, +q #�t      3    , +� #ߘ +d #ߘ +d %�t +� %�t +� #ߘ      3    , y4 %�� �� %�� �� 'T y4 'T y4 %��      3    , q@ 6< |� 6< |� �� q@ �� q@ 6<      3    , 4L 
�` @ 
�` @ � 4L � 4L 
�`      3    , q  �� |� �� |� ø q  ø q  ��      3    , Լ �� �t �� �t 7� Լ 7� Լ ��      3    , �@ 	�h �� 	�h �� 	׈ �@ 	׈ �@ 	�h      3    , �� � �� � �� �P �� �P �� �      3    ,  0< ��  ;� ��  ;� 0   0< 0   0< ��      3    , "�  �0 "l  �0 "l �� "� �� "�  �0      3    , !�� �� !�H �� !�H �0 !�� �0 !�� ��      3    , �h f< �  f< �  �l �h �l �h f<      3    , ]t �d i, �d i, � ]t � ]t �d      3    , �l #�� �$ #�� �$ #�� �l #�� �l #��      3    , �  @p � @p � :L �  :L �  @p      3    , � #�t �� #�t �� %� � %� � #�t      3    , �� #�t �x #�t �x $�< �� $�< �� #�t      3    , �� �, �l �, �l q� �� q� �� �,      3    , �� t �� t �� 6� �� 6� �� t      3    , op �| {( �| {( �� op �� op �|      3    , Z �| e� �| e� �� Z �� Z �|      3    , &� 
�P 2� 
�P 2� � &� � &� 
�P      3    , �� � �x � �x �� �� �� �� �      3    , �< �$ �� �$ �� :L �< :L �< �$      3    , KT !G� W !G� W !� KT !� KT !G�      3    , W0 "^� b� "^� b� #�� W0 #�� W0 "^�      3    , 9� !�� Ex !�� Ex "j� 9� "j� 9� !��      3    , 3� K0 ?P K0 ?P nX 3� nX 3� K0      3    , (�� #�� (� #�� (� #�� (�� #�� (�� #��      3    , 6< 	?0 A� 	?0 A� 	bX 6< 	bX 6< 	?0      3    , �0 K0 �� K0 �� nX �0 nX �0 K0      3    , � � �� � �� 7� � 7� � �      3    , �X %�L � %�L � %�t �X %�t �X %�L      3    , ]0 �� h� �� h� �T ]0 �T ]0 ��      3    , �p � ( � ( �� �p �� �p �      3    , �4 !�< �� !�< �� !�d �4 !�d �4 !�<      3    , �d !�� � !�� � "�� �d "�� �d !��      3    , � [| �< [| �< �� � �� � [|      3    , (�� � (� � (� vp (�� vp (�� �      3    , )�  � )�� � )�� C� )�  C� )�  �      3    , (� %�L (� %�L (� %�t (� %�t (� %�L      3    , %E %�L %P� %�L %P� %�� %E %�� %E %�L      3    , &�� d� &�� d� &�� �� &�� �� &�� d�      3    , �� �P h �P h ,� �� ,� �� �P      3    , �H �� �  �� �   �d �H  �d �H ��      3    , �   Ĭ ��  Ĭ �� !�d �  !�d �   Ĭ      3    , Y� � e@ � e@ y4 Y� y4 Y� �      3    , t � (, � (, 	� t 	� t �      3    , !P i� - i� - � !P � !P i�      3    , �� 	u� �| 	u� �| u� �� u� �� 	u�      3    , _$ !�< j� !�< j� !�d _$ !�d _$ !�<      3    , G� !�< SH !�< SH !�d G� !�d G� !�<      3    , M  � X� � X� =� M  =� M  �      3    , �� �  �  7� �� 7� �� �      3    , %�� �� %׀ �� %׀ �� %�� �� %�� ��      3    , �� �D � �D � �l �� �l �� �D      3    , !9� �� !E� �� !E�  � !9�  � !9� ��      3    , !� � !�\ � !�\ � !� � !� �      3    , 'e� � 'q� � 'q� 2� 'e� 2� 'e� �      3    , ,6\ � ,B � ,B 0  ,6\ 0  ,6\ �      3    , +o$ � +z� � +z� 0  +o$ 0  +o$ �      3    , 	{� �d 	�t �d 	�t �l 	{� �l 	{� �d      3    , *k` 	Ӡ *w 	Ӡ *w � *k` � *k` 	Ӡ      3    , �� � Ҁ � Ҁ V �� V �� �      3    , ;� � GH � GH �4 ;� �4 ;� �      3    ,   |� (� |� (� ��   ��   |�      3    , #CX �D #O �D #O �l #CX �l #CX �D      3    , a� 7� m8 7� m8 	bX a� 	bX a� 7�      3    , � 	j( %< 	j( %< 	�0 � 	�0 � 	j(      3    , &�� � &͘ � &͘ , &�� , &�� �      3    , �< � �� � �� �0 �< �0 �< �      3    , P t� ' t� ' 0  P 0  P t�      3    , H 	u� #  	u� #  	�0 H 	�0 H 	u�      3    , � K0 �� K0 �� �� � �� � K0      3    , �� 	u� �� 	u� �� 	� �� 	� �� 	u�      3    , �� K0 �8 K0 �8 	J� �� 	J� �� K0      3    , Լ � �t � �t )  Լ )  Լ �      3    , f� �� rd �� rd ø f� ø f� ��      3    , &Ǽ 
� &�t 
� &�t �� &Ǽ �� &Ǽ 
�      3    , (ul 	u� (�$ 	u� (�$ 
+� (ul 
+� (ul 	u�      3    , %� �d 1� �d 1� �T %� �T %� �d      3    , %� �` 1� �` 1� �l %� �l %� �`      3    , )�p � )�( � )�( 2� )�p 2� )�p �      3    , +� � +@ � +@ 2� +� 2� +� �      3    , 	�� � 	�P � 	�P �0 	�� �0 	�� �      3    , N� � Z@ � Z@ �0 N� �0 N� �      3    , �0 ʬ �� ʬ �� "�� �0 "�� �0 ʬ      3    , *�� z� *ڴ z� *ڴ :L *�� :L *�� z�      3    , | �� 4 �� 4 :L | :L | ��      3    , u � �� � �� �l u �l u �      3    , �| � �4 � �4 �l �| �l �| �      3    , �$ i� �� i� �� � �$ � �$ i�      3    , �� �  �H �  �H �P �� �P �� �       3    , Fl d� R$ d� R$ �� Fl �� Fl d�      3    , 	�H t� 	�  t� 	�  �� 	�H �� 	�H t�      3    , �\ � � � � � �\ � �\ �      3    , "� �� "� �� "� ø "� ø "� ��      3    , #� �� #�� �� #�� ø #� ø #� ��      3    , ې � �H � �H ,� ې ,� ې �      3    , )$ d� 4� d� 4� �� )$ �� )$ d�      3    , � "� �� "� �� #�( � #�( � "�      3    , �� �� а �� а ø �� ø �� ��      3    ,  A� �  M� �  M� )   A� )   A� �      3    , !, � !� � !� )  !, )  !, �      3    , �� M� �� M� �� j� �� j� �� M�      3    , Gl  �� S$  �� S$  ި Gl  ި Gl  ��      3    , O<  �0 Z�  �0 Z� [� O< [� O<  �0      3    , �H Z� �  Z� �  	bX �H 	bX �H Z�      3    , � � �� � �� �� � �� � �      3    , *X �d *% �d *% �� *X �� *X �d      3    , %� � %�� � %�� �� %� �� %� �      3    , +� d� +�� d� +�� �� +� �� +� d�      3    , -p d� -( d� -( �� -p �� -p d�      3    , �� ( �� ( �� 0  �� 0  �� (      3    , 	y� �� 	�� �� 	�� � 	y� � 	y� ��      3    , �X �� � �� � 	bX �X 	bX �X ��      3    , �� �� h �� h 	bX �� 	bX �� ��      3    , { "� �� "� �� #ݤ { #ݤ { "�      3    , (, �< 3� �< 3� !S@ (, !S@ (, �<      3    , �0 %�L �� %�L �� %�t �0 %�t �0 %�L      3    , � %�L �d %�L �d %�t � %�t � %�L      3    , �h 	� �  	� �  �0 �h �0 �h 	�      3    , v� i� �� i� �� � v� � v� i�      3    , g� i� s8 i� s8 � g� � g� i�      3    , �<  �x ��  �x �� [� �< [� �<  �x      3    , � 
�` �� 
�` �� � � � � 
�`      3    , %�`  �� %�  �� %�  ި %�`  ި %�`  ��      3    , �� �X � �X � 7� �� 7� �� �X      3    , �� �� �@ �� �@ 0  �� 0  �� ��      3    , )l �� 5$ �� 5$ �� )l �� )l ��      3    , �� =� � =� � a �� a �� =�      3    , � t� � t� � �� � �� � t�      3    , 4, �D ?� �D ?� �l 4, �l 4, �D      3    , ]� =� iP =� iP a ]� a ]� =�      3    ,  �, #�t  �� #�t  �� $�<  �, $�<  �, #�t      3    , F� %�� RH %�� RH &$ F� &$ F� %��      3    , �l !(H �$ !(H �$ !�d �l !�d �l !(H      3    , �0 $f\ � $f\ � %�t �0 %�t �0 $f\      3    , *�� 	j( *�� 	j( *�� 
� *�� 
� *�� 	j(      3    , &�� 
�P 'H 
�P 'H B@ &�� B@ &�� 
�P      3    , ,�� C� ,�h C� ,�h /H ,�� /H ,�� C�      3    , }� �� �@ �� �@ nT }� nT }� ��      3    , � 	u� �� 	u� �� 	� � 	� � 	u�      3    , � ?t �� ?t �� �� � �� � ?t      3    , x< �d �� �d �� K, x< K, x< �d      3    , �   d ��  d �� � �  � �   d      3    , ut !, �, !, �, B< ut B< ut !,      3    , l� K0 x` K0 x` fd l� fd l� K0      3    , "9� #ߘ "Ep #ߘ "Ep %� "9� %� "9� #ߘ      3    , �� K0 �� K0 �� �� �� �� �� K0      3    , �� ^� �` ^� �` �� �� �� �� ^�      3    , �� � �� � �� "� �� "� �� �      3    , X� �� dH �� dH �� X� �� X� ��      3    , �� x �L x �L #  �� #  �� x      3    , s\ 	u�  	u�  '0 s\ '0 s\ 	u�      3    , v� �� �h �� �h x v� x v� ��      3    , !f� �� !r� �� !r�  !f�  !f� ��      3    , !f� �P !r� �P !r� �l !f� �l !f� �P      3    , � M� �� M� �� (� � (� � M�      3    , 
j C� 
u� C� 
u� �� 
j �� 
j C�      3    , f� |� r� |� r� �� f� �� f� |�      3    , �� J �� J �� �D �� �D �� J      3    , ,�p h ,�( h ,�( 	bX ,�p 	bX ,�p h      3    , -�� ld -�� ld -�� 8 -�� 8 -�� ld      3    , �� J �� J �� �\ �� �\ �� J      3    , �t _D �, _D �, �T �t �T �t _D      3    , _� M� k� M� k� j� _� j� _� M�      3    , �� �< �� �< �� �d �� �d �� �<      3    , +�p |� +�( |� +�( �� +�p �� +�p |�      3    , \� �l h� �l h� a \� a \� �l      3    , �� L �h L �h �l �� �l �� L      3    , X� eD dp eD dp �� X� �� X� eD      3    , �� 	� �� 	� �� �0 �� �0 �� 	�      3    , �H �d �  �d �  �� �H �� �H �d      3    , �@ � �� � �� �� �@ �� �@ �      3    , H� �, T` �, T` � H� � H� �,      3    , 
�P !�� 
� !�� 
� " 
�P " 
�P !��      3    , )�� �< )�� �< )��  �d )��  �d )�� �<      3    , (PP �� (\ �� (\ �d (PP �d (PP ��      3    , |� t� �H t� �H �| |� �| |� t�      3    , � ET �� ET �� C< � C< � ET      3    , b \ m� \ m� 	bX b 	bX b \      3    , 	�� �� 	�8 �� 	�8 0  	�� 0  	�� ��      3    , wD 4 �� 4 �� �� wD �� wD 4      3    , $� =� 0� =� 0� a $� a $� =�      3    , �� K0 �< K0 �< Z� �� Z� �� K0      3    , �� M�  M�  I� �� I� �� M�      3    , ( =� � =� � a ( a ( =�      3    , � �X � �X � 7� � 7� � �X      3    , tx �X �0 �X �0 7� tx 7� tx �X      3    , �� b� � b� � 	bX �� 	bX �� b�      3    , )� � 5h � 5h 0  )� 0  )� �      3    , )�p M� )�( M� )�( p� )�p p� )�p M�      3    , � |� � |� � �� � �� � |�      3    , 	� �� x �� x 3, 	� 3, 	� ��      3    , � � �� � �� �4 � �4 � �      3    , 5   �0 @�  �0 @� X 5  X 5   �0      3    , Ll  �0 X$  �0 X$ X Ll X Ll  �0      3    ,  
�h � 
�h � ��  ��  
�h      3    , �L 	u� � 	u� � 
�  �L 
�  �L 	u�      3    , &� �0 2\ �0 2\ C` &� C` &� �0      3    , �P  �0 �  �0 � ~� �P ~� �P  �0      3    , 
� � 
)� � 
)� � 
� � 
� �      3    , 
!� � 
-x � 
-x B@ 
!� B@ 
!� �      3    , �\ C� � C� � f� �\ f� �\ C�      3    , �� [ Ƥ [ Ƥ �H �� �H �� [      3    , �� !`� �� !`� �� !� �� !� �� !`�      3    , .P %�� : %�� : &$ .P &$ .P %��      3    , dH � p  � p  �� dH �� dH �      3    , D �� (� �� (� YH D YH D ��      3    , e� M� q@ M� q@ 0  e� 0  e� M�      3    , "�� �\ "� �\ "� �� "�� �� "�� �\      3    , #)� K0 #5� K0 #5� 	J� #)� 	J� #)� K0      3    , 	�� K0 	�� K0 	�� 	bX 	�� 	bX 	�� K0      3    , �� 	u�  8 	u�  8 	� �� 	� �� 	u�      3    , �| 	?0 �4 	?0 �4 	bX �| 	bX �| 	?0      3    , x� G� �` G� �` E� x� E� x� G�      3    , U\ t� a t� a �� U\ �� U\ t�      3    , !� � !�P � !�P <d !� <d !� �      3    , 
h #�t 
s� #�t 
s� %�� 
h %�� 
h #�t      3    , *�, �, *�� �, *�� H� *�, H� *�, �,      3    , )� !�< )| !�< )| !�d )� !�d )� !�<      3    , l� %�L x� %�L x� %�t l� %�t l� %�L      3    , |l %�L �$ %�L �$ %�P |l %�P |l %�L      3    , Z� C� f� C� f� f� Z� f� Z� C�      3    , ^H ~@ j  ~@ j  7� ^H 7� ^H ~@      3    , �� � �8 � �8 �4 �� �4 �� �      3    , 
�t �� 
, �� 
, � 
�t � 
�t ��      3    , � ~� �` ~� �` �d � �d � ~�      3    , �4 %�L �� %�L �� %�t �4 %�t �4 %�L      3    , @ ,� K� ,� K� � @ � @ ,�      3    , ~� �� �@ �� �@ � ~� � ~� ��      3    , 
� � 
�� � 
�� _� 
� _� 
� �      3    , ,\ 	?0 8 	?0 8 	bX ,\ 	bX ,\ 	?0      3    , W� 7� c� 7� c� 	bX W� 	bX W� 7�      3    , � �� x �� x qh � qh � ��      3    , �� =� � =� � f� �� f� �� =�      3    , :l F� F$ F� F$ � :l � :l F�      3    , !� i� -t i� -t � !� � !� i�      3    , +q �d +|� �d +|� C\ +q C\ +q �d      3    , ,@ � ,� � ,�  ,@  ,@ �      3    , �� �� �\ �� �\ �� �� �� �� ��      3    , hT �( t �( t �$ hT �$ hT �(      3    , .� $ � .� $ � .� $+� .� $+� .� $ �      3    , )�� #�t )� #�t )� $� )�� $� )�� #�t      3    , �d %�D � %�D � 'T �d 'T �d %�D      3    , rd %�� ~ %�� ~ &$ rd &$ rd %��      3    , �� C� �x C� �x f� �� f� �� C�      3    , 7� d� C� d� C� �� 7� �� 7� d�      3    , �$ �� �� �� �� � �$ � �$ ��      3    , (� �L 4� �L 4� I� (� I� (� �L      3    , 
�4 M� 
�� M� 
�� p� 
�4 p� 
�4 M�      3    , "5� �| "A� �| "A� �� "5� �� "5� �|      3    , #�� �| #�d �| #�d �� #�� �� #�� �|      3    , �H t� �  t� �  �� �H �� �H t�      3    , $�| �, $�4 �, $�4 �T $�| �T $�| �,      3    , &-p �, &9( �, &9( �T &-p �T &-p �,      3    , � �$ *� �$ *� �� � �� � �$      3    , �l �d �$ �d �$ � �l � �l �d      3    , �� �� �d �� �d �4 �� �4 �� ��      3    , �0 f< �� f< �� �l �0 �l �0 f<      3    , .G� d� .S` d� .S` �� .G� �� .G� d�      3    , -�P d� -� d� -� �� -�P �� -�P d�      3    ,  �� �|  �� �|  �� ��  �� ��  �� �|      3    , ֈ �| �@ �| �@ � ֈ � ֈ �|      3    , )� i� )� i� )� � )� � )� i�      3    , )� �� )� �� )� < )� < )� ��      3    , -p� #ټ -|� #ټ -|� $� -p� $� -p� #ټ      3    , .� #�t .� #�t .� $� .� $� .� #�t      3    , �� �| �� �| �� �� �� �� �� �|      3    , ' �� 2� �� 2� )  ' )  ' ��      3    , ¼ �� �t �� �t c0 ¼ c0 ¼ ��      3    , (�� �� (�h �� (�h ø (�� ø (�� ��      3    , -� !�� 9P !�� 9P " -� " -� !��      3    , | �� 4 �� 4 �� | �� | ��      3    , � �� �� �� �� Rl � Rl � ��      3    , ?� M� Kt M� Kt j� ?� j� ?� M�      3    , 2 �� =� �� =� �� 2 �� 2 ��      3    , Đ � �H � �H 6� Đ 6� Đ �      3    , 	�� 	u� 	�8 	u� 	�8 \ 	�� \ 	�� 	u�      3    , v�  d ��  d �� �4 v� �4 v�  d      3    , 
� �, t �, t �T 
� �T 
� �,      3    , P %�L ! %�L ! %�t P %�t P %�L      3    , "�P �4 "� �4 "� <` "�P <` "�P �4      3    , (g� d� (sx d� (sx �� (g� �� (g� d�      3    , *@ �� *(� �� *(� � *@ � *@ ��      3    , *@h ( *L  ( *L  0  *@h 0  *@h (      3    , %y� t� %�x t� %�x �� %y� �� %y� t�      3    , �� �� ̠ �� ̠ �� �� �� �� ��      3    , �\ �, � �, � �4 �\ �4 �\ �,      3    , �� � �� � �� �0 �� �0 �� �      3    , �  � �� � �� �0 �  �0 �  �      3    , �� 	u� �� 	u� �� 	� �� 	� �� 	u�      3    , +� 
d( 7� 
d( 7� � +� � +� 
d(      3    , �� �@ �| �@ �| � �� � �� �@      3    , � �� )h �� )h �\ � �\ � ��      3    , g� $�� s� $�� s� %�@ g� %�@ g� $��      3    , � #�t h #�t h %� � %� � #�t      3    , M$ �< X� �< X� !0 M$ !0 M$ �<      3    , 4� C� @� C� @� f� 4� f� 4� C�      3    , � �� x �� x �� � �� � ��      3    , �d �d � �d � � �d � �d �d      3    , ^l C� j$ C� j$ �� ^l �� ^l C�      3    , �p K0 �( K0 �( nX �p nX �p K0      3    , 	�p �, 	�( �, 	�( �T 	�p �T 	�p �,      3    , e� f< qh f< qh �l e� �l e� f<      3    , � M� l M� l � � � � M�      3    , �� M� �@ M� �@ � �� � �� M�      3    , $�� M� $�� M� $�� �$ $�� �$ $�� M�      3    , *�P �` *� �` *� nX *�P nX *�P �`      3    , %#� K0 %/� K0 %/� nX %#� nX %#� K0      3    , 6� �� Bd �� Bd  6�  6� ��      3    , � L � L � �4 � �4 � L      3    , � �( �� �( �� �P � �P � �(      3    , (� t� (�� t� (�� �� (� �� (� t�      3    , )�h t� )�  t� )�  �� )�h �� )�h t�      3    , 0   �� ;�  �� ;�  ި 0   ި 0   ��      3    , ]� 	u� iP 	u� iP 	�X ]� 	�X ]� 	u�      3    , x� �  �� �  �� �P x� �P x� �       3    , +4 i� +$� i� +$� � +4 � +4 i�      3    , )JP $ )V $ )V :L )JP :L )JP $      3    , !�P 	u� " 	u� " 
h !�P 
h !�P 	u�      3    , � !�< �� !�< �� !�d � !�d � !�<      3    , �� �< �@ �< �@  �d ��  �d �� �<      3    , %� !�L 18 !�L 18 " %� " %� !�L      3    , �� � �| � �| � �� � �� �      3    , �D � �� � �� ,� �D ,� �D �      3    , �0 ', �� ', �� 6� �0 6� �0 ',      3    , �@ � �� � �� 2� �@ 2� �@ �      3    , 'i� M� 'u� M� 'u� �� 'i� �� 'i� M�      3    , �� �, Ҥ �, Ҥ � �� � �� �,      3    , E� M� Qt M� Qt p� E� p� E� M�      3    , U� �, a\ �, a\ N� U� N� U� �,      3    , �� C ؤ C ؤ �l �� �l �� C      3    , �� B �8 B �8 �\ �� �\ �� B      3    , /� =� ;� =� ;� a /� a /� =�      3    , #� �( #�� �( #�� �P #� �P #� �(      3    , )  	?0 )� 	?0 )� 	bX )  	bX )  	?0      3    , �\ 	p � 	p � 
H� �\ 
H� �\ 	p      3    , m� 
= y� 
= y� �� m� �� m� 
=      3    , ݈ 	�x �@ 	�x �@ �� ݈ �� ݈ 	�x      3    , k� �� wh �� wh a k� a k� ��      3    , � %�� � %�� � &$ � &$ � %��      3    ,  � %�� ,8 %�� ,8 &$  � &$  � %��      3    , pL !Kp | !Kp | #ݤ pL #ݤ pL !Kp      3    , 	4 � � � � 0  	4 0  	4 �      3    , �� � � � � 0  �� 0  �� �      3    , �� e� �x e� �x � �� � �� e�      3    , �� �� �H �� �H �p �� �p �� ��      3    , "�T M� "� M� "� �L "�T �L "�T M�      3    ,  � #��  � #��  � #��  � #��  � #��      3    , &�� � &ˤ � &ˤ 7� &�� 7� &�� �      3    , #
� 	u� #l 	u� #l 	�0 #
� 	�0 #
� 	u�      3    , �� �, x �, x �T �� �T �� �,      3    , 
1` J 
= J 
= �T 
1` �T 
1` J      3    , e@ #�� p� #�� p� #�� e@ #�� e@ #��      3    , J0 #�� U� #�� U� #�� J0 #�� J0 #��      3    , #�� �� #�x �� #�x � #�� � #�� ��      3    ,  � �  �� �  �� �0  � �0  � �      3    , |� hT �h hT �h �l |� �l |� hT      3    , "7� =� "C| =� "C| �  "7� �  "7� =�   	   3    !    �  '7 � '7 �      3    , �� �� �d �� �d � �� � �� ��      3    , @ �8 )� �8 )� )  @ )  @ �8      3    , $0 � $%� � $%� )  $0 )  $0 �      3    , %�� M� &x M� &x �$ %�� �$ %�� M�      3    , *�  �T *L  �T *L �� *� �� *�  �T      3    , � �� �� �� �� 0  � 0  � ��      3    , +Q� L +]� L +]� f� +Q� f� +Q� L      3    , �� !� �� !� �� !�d �� !�d �� !�      3    , &�$ �� &�� �� &�� 	bX &�$ 	bX &�$ ��      3    , '!� �� '-L �� '-L 	�X '!� 	�X '!� ��      3    , ۴ �, �l �, �l �T ۴ �T ۴ �,      3    , c, �< n� �< n� �� c, �� c, �<      3    , .P t� : t� : �� .P �� .P t�      3    , -A� �, -M� �, -M� �t -A� �t -A� �,      3    , ̤ :l �\ :l �\ m4 ̤ m4 ̤ :l      3    , Q� �, ]T �, ]T �T Q� �T Q� �,      3    ,  Qp 
ɸ  ]( 
ɸ  ]( �  Qp �  Qp 
ɸ      3    , #�� 	u� $� 	u� $� 	� #�� 	� #�� 	u�      3    , �� � �d � �d �� �� �� �� �      3    , AD �4 L� �4 L� 6� AD 6� AD �4      3    , %/� =� %;@ =� %;@ a %/� a %/� =�      3    , %�� =� %Ә =� %Ә a %�� a %�� =�      3    , %` �� 1 �� 1 c0 %` c0 %` ��      3    , �  t� �� t� �� �� �  �� �  t�      3    , � � �� � �� )  � )  � �      3    , *�@ C� *�� C� *�� �� *�@ �� *�@ C�      3    , *�X U` *� U` *� 0  *�X 0  *�X U`      3    , #�� � $
� � $
� 0  #�� 0  #�� �      3    , +�� �� +�h �� +�h ø +�� ø +�� ��      3    , �< !�� �� !�� �� " �< " �< !��      3    , �� !�� � !�� � " �� " �� !��      3    , �( � �� � �� )  �( )  �( �      3    , i0 �� t� �� t� �� i0 �� i0 ��      3    , � � �� � �� �0 � �0 � �      3    , 
�P � 
� � 
� �4 
�P �4 
�P �      3    , � }� �H }� �H 
�  � 
�  � }�      3    , S� �� _d �� _d �� S� �� S� ��   	   3    !    �P  �� 4t �� &x +  ,VR_LEFT_VERTICAL_BUS      3    , *�� .P *�P .P *�P 5� *�� 5� *�� .P      3    , ![ �( !f� �( !f� �P ![ �P ![ �(      3    , *6� 	?0 *B\ 	?0 *B\ 	bX *6� 	bX *6� 	?0      3    , '0 � 2� � 2� �0 '0 �0 '0 �      3    , 	Ѭ !�< 	�d !�< 	�d !�d 	Ѭ !�d 	Ѭ !�<      3    , �� �D Θ �D Θ �l �� �l �� �D      3    , �� �D ̀ �D ̀ �l �� �l �� �D      3    , �x !�� �0 !�� �0 $� �x $� �x !��      3    , �< K0 �� K0 �� f� �< f� �< K0      3    , �L Z� � Z� � 	bX �L 	bX �L Z�      3    , Z� M� f� M� f� p� Z� p� Z� M�      3    , f� M� r� M� r� p� f� p� f� M�      3    , +�� 	p +�x 	p +�x � +�� � +�� 	p      3    , +]� K0 +iH K0 +iH hX +]� hX +]� K0      3    , ې t� �H t� �H l� ې l� ې t�      3    , 	0 �� � �� �  	0  	0 ��      3    , � #�t � #�t � $+� � $+� � #�t      3    , !n� !�< !zP !�< !zP !�d !n� !�d !n� !�<      3    , #5� � #Ad � #Ad 0  #5� 0  #5� �      3    , 80 x� C� x� C� �� 80 �� 80 x�      3    , �� � �x � �x �t �� �t �� �      3    , �� �� �� �� �� 6� �� 6� �� ��      3    , � h� � h� � (L � (L � h�      3    , V� n� bT n� bT �� V� �� V� n�      3    , 1� \ =� \ =� 	bX 1� 	bX 1� \      3    , �� #�t d #�t d $�d �� $�d �� #�t      3    , �| �  �4 �  �4 <d �| <d �| �       3    , �| �� �4 �� �4 0  �| 0  �| ��      3    , )�� %�t )�� %�t )�� &= )�� &= )�� %�t      3    , 'T\  �0 '`  �0 '` $� 'T\ $� 'T\  �0      3    , (�l  �0 (�$  �0 (�$ $� (�l $� (�l  �0      3    , (�x @ (�0 @ (�0 �� (�x �� (�x @      3    , /H �$ ;  �$ ;  :L /H :L /H �$      3    , :� $�� FH $�� FH %�P :� %�P :� $��      3    , | � �4 � �4 �0 | �0 | �      3    , 
H� S� 
T� S� 
T� �0 
H� �0 
H� S�      3    , 
H� �� 
T� �� 
T� �� 
H� �� 
H� ��      3    , � "l d "l d #�� � #�� � "l      3    ,  � %�$ ,| %�$ ,| %�t  � %�t  � %�$      3    , � � � � � )  � )  � �      3    , & H 1� H 1� �4 & �4 & H      3    , �� C� h C� h f� �� f� �� C�      3    , 4� � @H � @H �0 4� �0 4� �      3    , $ � � � � �� $ �� $ �      3    , � a� � a� � �P � �P � a�      3    , � �( �� �( �� �P � �P � �(      3    , 1� �( =� �( =� F 1� F 1� �(      3    , "b� �, "nt �, "nt k� "b� k� "b� �,      3    , )�p �d )�( �d )�( Ah )�p Ah )�p �d      3    ,   t� � t� � �   �   t�      3    , �� � h � h 0  �� 0  �� �      3    , }� $ �d $ �d :L }� :L }� $      3    , �| �� �4 �� �4 !�d �| !�d �| ��      3    , �� �< �l �< �l !0 �� !0 �� �<      3    , �h #�� �  #�� �  $r �h $r �h #��      3    , �� $ Ƥ $ Ƥ :L �� :L �� $      3    , �0 p$ � p$ � �l �0 �l �0 p$      3    , � d� �� d� �� �� � �� � d�      3    , 9� |� EP |� EP �� 9� �� 9� |�      3    , N� |� Z� |� Z� �� N� �� N� |�      3    , #�� 
�P $� 
�P $� :L #�� :L #�� 
�P      3    , 	P =�  =�  a 	P a 	P =�      3    , 0� C� <@ C� <@ �� 0� �� 0� C�      3    , 
5H � 
A  � 
A  7� 
5H 7� 
5H �      3    , �� $ ɐ $ ɐ :L �� :L �� $      3    , '#�  �0 '/@  �0 '/@ kH '#� kH '#�  �0      3    , *@ =� 5� =� 5� GH *@ GH *@ =�      3    , .( � 9� � 9� 5� .( 5� .( �      3    , � %�L #� %�L #� %�t � %�t � %�L      3    , �0 � �� � �� �4 �0 �4 �0 �      3    , �� �� 	� �� 	� �� �� �� �� ��      3    , Y� C� e@ C� e@ �  Y� �  Y� C�      3    , 6` �h B �h B Z� 6` Z� 6` �h      3    , Z� ^� f� ^� f� 	bX Z� 	bX Z� ^�      3    , � �� �< �� �< �� � �� � ��      3    , �� !�� �x !�� �x #�| �� #�| �� !��      3    , Ð #�t �H #�t �H $� Ð $� Ð #�t      3    , -�� \ -�h \ -�h 6� -�� 6� -�� \      3    , � =� �� =� �� a � a � =�      3    , x` �� � �� � �� x` �� x` ��      3    , < \ $� \ $� B< < B< < \      3    , %< �4 0� �4 0� 6� %< 6� %< �4      3    , �� %�L �d %�L �d %�t �� %�t �� %�L      3    , �� %�L �\ %�L �\ %�t �� %�t �� %�L      3    , �� �d � �d � �� �� �� �� �d      3    , *,� �D *8� �D *8� �l *,� �l *,� �D      3    , +m0 �D +x� �D +x� �l +m0 �l +m0 �D      3    , � %�\ �� %�\ �� &3L � &3L � %�\      3    , )2� �| )>� �| )>� �� )2� �� )2� �|      3    , " T � ", � ", y4 " T y4 " T �      3    , -X C� - C� - �� -X �� -X C�      3    , -�l F� -�$ F� -�$ �4 -�l �4 -�l F�      3    , $P� 
�x $\� 
�x $\� � $P� � $P� 
�x      3    , � $ �� $ �� :L � :L � $      3    , �� C� �� C� �� �� �� �� �� C�      3    , ( a| � a| � g4 ( g4 ( a|      3    , (P J 4 J 4 g4 (P g4 (P J      3    , Ѩ �( �` �( �` �P Ѩ �P Ѩ �(      3    , 	�H �4 	�  �4 	�  �� 	�H �� 	�H �4      3    , 	/� ET 	;H ET 	;H nX 	/� nX 	/� ET      3    , )>� $jD )JP $jD )JP %�� )>� %�� )>� $jD      3    , �d "�� � "�� � #�� �d #�� �d "��      3    , .&t �� .2, �� .2, Xl .&t Xl .&t ��      3    , Ml �, Y$ �, Y$ �T Ml �T Ml �,      3    , k� �� w� �� w� �� k� �� k� ��      3    , @� M� L� M� L� �� @� �� @� M�      3    , "d� 	 "ph 	 "ph 	bX "d� 	bX "d� 	      3    , (PP � (\ � (\ 	n (PP 	n (PP �      3    , � d� �� d� �� �� � �� � d�      3    , � \ �� \ �� 6� � 6� � \      3    , (B� F� (N\ F� (N\ � (B� � (B� F�      3    , �P d� � d� � �� �P �� �P d�      3    , �P d� � d� � �� �P �� �P d�      3    , 24 � =� � =� �� 24 �� 24 �      3    , t� _D �T _D �T a t� a t� _D      3    , �` � � � � )  �` )  �` �      3    , #� � /� � /� �0 #� �0 #� �      3    , �� � 	� � 	� �0 �� �0 �� �      3    , �� � � � � 0  �� 0  �� �      3    , �p �h �( �h �( K0 �p K0 �p �h      3    , Z� �| fd �| fd �� Z� �� Z� �|      3    , �< 	?0 �� 	?0 �� 	bX �< 	bX �< 	?0      3    , 
�� �d 
�x �d 
�x ( 
�� ( 
�� �d      3    , Ԙ 	u� �P 	u� �P 	� Ԙ 	� Ԙ 	u�      3    , �� *h �L *h �L 0  �� 0  �� *h      3    , k� 	u� w� 	u� w� 	� k� 	� k� 	u�      3    , 6<  �0 A�  �0 A� X 6< X 6<  �0      3    , !��  �0 !�  �0 !� X !�� X !��  �0      3    , �� �� �� �� �� 4 �� 4 �� ��      3    , 
� h� L h� L nT 
� nT 
� h�      3    , Mh �4 Y  �4 Y  B< Mh B< Mh �4      3    , �� #� А #� А �l �� �l �� #�      3    , ,� �d 88 �d 88 �� ,� �� ,� �d      3    , � J @ J @ g4 � g4 � J      3    , � � *d � *d F$ � F$ � �      3    , � 	u� �� 	u� �� 	�0 � 	�0 � 	u�      3    , �0 	?0 �� 	?0 �� 	bX �0 	bX �0 	?0      3    , �� �, �H �, �H �T �� �T �� �,      3    , �� J �� J �� m4 �� m4 �� J      3    , "� t� #� t� #� � "� � "� t�      3    , �� �� �� �� �� �� �� �� �� ��      3    , �l �, �$ �, �$ | �l | �l �,      3    , 	T� !Kp 	`d !Kp 	`d !�d 	T� !�d 	T� !Kp      3    , �� �< �� �< �� !W( �� !W( �� �<      3    , ,g0 �l ,r� �l ,r� a ,g0 a ,g0 �l      3    , �� M� �l M� �l �$ �� �$ �� M�      3    , �� = � = � �l �� �l �� =      3    , *0� |� *<� |� *<� �� *0� �� *0� |�      3    , �l �( �$ �( �$ �P �l �P �l �(      3    , s� �( 8 �( 8 �P s� �P s� �(      3    , 
  � 
� � 
� 7� 
  7� 
  �      3    , Ŭ C� �d C� �d f� Ŭ f� Ŭ C�      3    , � �� � �� � 0  � 0  � ��      3    , 5� s A� s A� �� 5� �� 5� s      3    , W� v� cP v� cP �D W� �D W� v�      3    , *� C� 6� C� 6� f� *� f� *� C�   	   3    !    �  �4 Q �4 T�      3    , � ,� �` ,� �` �0 � �0 � ,�      3    , � �� �` �� �` ?� � ?� � ��      3    , %q� J %}� J %}� m4 %q� m4 %q� J      3    ,  �P $ !	 $ !	 p�  �P p�  �P $      3    , $0 �d $%� �d $%� �L $0 �L $0 �d      3    , 2\ �, > �, > /� 2\ /� 2\ �,      3    , !zP � !� � !� 7� !zP 7� !zP �      3    , !�0 
d( !�� 
d( !�� � !�0 � !�0 
d(      3    , %)� �, %5d �, %5d | %)� | %)� �,      3    , ~d � � � � =� ~d =� ~d �      3    , F� 
= Rp 
= Rp �� F� �� F� 
=      3    , T` �� ` �� ` �� T` �� T` ��   	   3    !    �P  /=� 4t /=� &x +  ,VR_RIGHT_VERTICAL_BUS       3    , �0 �� �� �� ��  � �0  � �0 ��      3    , �D !�� �� !�� �� " �D " �D !��      3    , ְ �< �h �< �h �d ְ �d ְ �<      3    ,  � 7�  *` 7�  *` 	h4  � 	h4  � 7�      3    , )6� m| )B� m| )B� 6� )6� 6� )6� m|      3    , (m� $ (yT $ (yT :L (m� :L (m� $      3    , '� M� '�� M� '�� �t '� �t '� M�      3    , � M� �` M� �` p� � p� � M�      3    , J| � V4 � V4 F J| F J| �      3    , +�X C� +� C� +� _  +�X _  +�X C�      3    , *gx SH *s0 SH *s0 7� *gx 7� *gx SH      3    , ̀ #�t �8 #�t �8 $� ̀ $� ̀ #�t      3    , $d #�� 0 #�� 0 #�� $d #�� $d #��      3    , ƀ !�� �8 !�� �8 "�� ƀ "�� ƀ !��      3    , +q #�� +|� #�� +|� #�� +q #�� +q #��      3    , �� �� ˨ �� ˨ a �� a �� ��      3    , �� !$` Ô !$` Ô !� �� !� �� !$`      3    , � |� � |� � �� � �� � |�      3    , *[� �( *gx �( *gx �P *[� �P *[� �(      3    , (�� M� (� M� (� p� (�� p� (�� M�      3    , ,$� $ ,0� $ ,0� :L ,$� :L ,$� $      3    , ,G� t� ,S� t� ,S� �� ,G� �� ,G� t�      3    , � t� �@ t� �@ n� � n� � t�      3    , o, %�L z� %�L z� %�t o, %�t o, %�L      3    , K, %�� V� %�� V� &3L K, &3L K, %��      3    , z| �� �4 �� �4 �� z| �� z| ��      3    , $dh �( $p  �( $p  �P $dh �P $dh �(      3    , a| #�� m4 #�� m4 #�� a| #�� a| #��      3    , �p �< �( �< �(  �x �p  �x �p �<      3    , ]t #�� i, #�� i, #�� ]t #�� ]t #��      3    , wh i� �  i� �  � wh � wh i�      3    , �d 	f@  	f@  �� �d �� �d 	f@      3    , �\ � � � � 0  �\ 0  �\ �      3    , (� #�t (�� #�t (�� $x (� $x (� #�t      3    , '�X $� '� $� '� %�t '�X %�t '�X $�      3    , .p =� :( =� :( a .p a .p =�      3    , �� =� �@ =� �@ a �� a �� =�      3    , �$ A� �� A� �� �� �$ �� �$ A�      3    , �\ t� � t� � MD �\ MD �\ t�      3    , )a� � )mx � )mx �0 )a� �0 )a� �      3    , )�0 d� *� d� *� �� )�0 �� )�0 d�      3    , � �< �� �< �� !�� � !�� � �<      3    , �d !�< � !�< � !�d �d !�d �d !�<      3    , �$ !�� �� !�� �� "$< �$ "$< �$ !��      3    , $I M� $T� M� $T� �t $I �t $I M�      3    , "�� d� "�X d� "�X �� "�� �� "�� d�      3    , LH �D X  �D X  �H LH �H LH �D      3    , �0 �  �� �  �� �P �0 �P �0 �       3    , q� �� }@ �� }@ �� q� �� q� ��      3    , #K( t� #V� t� #V� pl #K( pl #K( t�      3    , &d  ?t &o� ?t &o� �� &d  �� &d  ?t      3    , g� %�� s� %�� s� &$ g� &$ g� %��      3    , 2| �� >4 �� >4 | 2| | 2| ��      3    , �`  �� �  �� �  ި �`  ި �`  ��      3    , 4  �� �  �� �  ި 4  ި 4  ��      3    , ` � k� � k� 0  ` 0  ` �      3    , 2X  �0 >  �0 > �� 2X �� 2X  �0      3    , ''p ";� '3( ";� '3( #�� ''p #�� ''p ";�      3    , #�, !�� #�� !�� #�� "Gd #�, "Gd #�, !��      3    , !�p �� !�( �� !�( �4 !�p �4 !�p ��      3    , !C� �< !OX �< !OX �� !C� �� !C� �<      3    , +m0 �( +x� �( +x� �P +m0 �P +m0 �(      3    , ,|� �( ,�d �( ,�d �P ,|� �P ,|� �(      3    , �� "�� �H "�� �H #�� �� #�� �� "��      3    , �� �� �� �� ��  ��  �� ��      3    , � #�t *� #�t *� $�L � $�L � #�t      3    , 6  �| A� �| A� �� 6  �� 6  �|      3    , %R� �� %^h �� %^h � %R� � %R� ��      3    , )�� �� )�� �� )�� � )�� � )�� ��      3    , %�� K0 %�� K0 %�� �� %�� �� %�� K0      3    , *��  �� *ڴ  �� *ڴ  ި *��  ި *��  ��      3    , )�T  �� )�  �� )�  ި )�T  ި )�T  ��      3    , � W0 �H W0 �H C` � C` � W0      3    , �l � �$ � �$ 0  �l 0  �l �      3    , �X �| � �| � a �X a �X �|      3    , �� M� �x M� �x �$ �� �$ �� M�      3    , $� �� $�� �� $�� a $� a $� ��      3    , 
�| J 
�4 J 
�4 �T 
�| �T 
�| J      3    , 
�� �� 8 �� 8 , 
�� , 
�� ��      3    , {� � �L � �L )  {� )  {� �      3    , :H n� F  n� F  �� :H �� :H n�      3    , "�` J "� J "� �l "�` �l "�` J      3    , %
l � %$ � %$ V %
l V %
l �      3    ,  0< ��  ;� ��  ;�   0<   0< ��      3    , U| � a4 � a4 �4 U| �4 U| �      3    , !  =� !� =� !� f� !  f� !  =�      3    , "h�  �� "tP  �� "tP  ި "h�  ި "h�  ��      3    , #/�  �� #;�  �� #;�  ި #/�  ި #/�  ��      3    , )�  � )��  � )�� kH )� kH )�  �      3    , ۴ "�D �l "�D �l #�� ۴ #�� ۴ "�D      3    , ��  ' 	
t  ' 	
t  ި ��  ި ��  '      3    , 	bX 	u� 	n 	u� 	n %� 	bX %� 	bX 	u�      3    , PX 	?0 \ 	?0 \ 	bX PX 	bX PX 	?0      3    , � $ �H $ �H :L � :L � $      3    , \ � % � % �0 \ �0 \ �      3    , �� �� �� �� ��  ��  �� ��      3    , :l !�< F$ !�< F$ !�d :l !�d :l !�<      3    , (�� J (�� J (�� �\ (�� �\ (�� J      3    , (ul �< (�$ �< (�$ �� (ul �� (ul �<      3    , ,�� � ,Ԑ � ,Ԑ 7� ,�� 7� ,�� �      3    , -�� h .@ h .@ 	bX -�� 	bX -�� h      3    , 	'� �� 	3x �� 	3x  	'�  	'� ��      3    , 
Zd �� 
f �� 
f  
Zd  
Zd ��      3    , V4 �� a� �� a�  V4  V4 ��      3    , �$ �  �� �  ��  �$  �$ �       3    , �� � Đ � Đ �P �� �P �� �      3    , �� �� �h �� �h �0 �� �0 �� ��      3    , . K0 .� K0 .� x . x . K0      3    , $p  !�� ${� !�� ${� " $p  " $p  !��      3    , P i� ! i� ! � P � P i�      3    , �� � �` � �` �� �� �� �� �      3    , � 28 L 28 L ;� � ;� � 28      3    , "�� � "�� � "�� #  "�� #  "�� �      3    , q� !�� }� !�� }� " q� " q� !��      3    , �  �0 	�  �0 	� <h � <h �  �0      3    , +(� �4 +4� �4 +4� �� +(� �� +(� �4      3    , w !�< �� !�< �� !�d w !�d w !�<      3    , �, #�� 	� #�� 	� #�� �, #�� �, #��      3    , $�X %�� $� %�� $� 'L� $�X 'L� $�X %��      3    , e� t� qD t� qD $ e� $ e� t�      3    , �P �4 � �4 � 6� �P 6� �P �4      3    , �L �� � �� � � �L � �L ��      3    , �� 
�P �d 
�P �d � �� � �� 
�P      3    , � �� �� �� �� �� � �� � ��      3    , �� 	u� �d 	u� �d 
H� �� 
H� �� 	u�      3    , %R� "^� %^h "^� %^h #�� %R� #�� %R� "^�      3    , 4p �$ @( �$ @( :L 4p :L 4p �$      3    , #?p �� #K( �� #K( @ #?p @ #?p ��      3    , + �h 6� �h 6� �4 + �4 + �h      3    , .zp � .�( � .�( 2� .zp 2� .zp �      3    , 	\| !�� 	h4 !�� 	h4 " 	\| " 	\| !��      3    , �< �� �� �� �� �� �< �� �< ��      3    , %�� �� %�@ �� %�@ �P %�� �P %�� ��      3    , �� � �� � �� �0 �� �0 �� �      3    , � �� �h �� �h  �  � ��      3    , �� M� �< M� �< l �� l �� M�      3    , 9� �l EP �l EP �\ 9� �\ 9� �l      3    , *@ 	 *(� 	 *(� 0  *@ 0  *@ 	      3    , +� %�� 7� %�� 7� &$ +� &$ +� %��      3    , � H �� H �� :L � :L � H      3    , )+ 	u� )6� 	u� )6� 	�0 )+ 	�0 )+ 	u�      3    , *�� 	u� +� 	u� +� 	�0 *�� 	�0 *�� 	u�      3    , #� C� #T C� #T f� #� f� #� C�      3    , 	 � � � � �0 	 �0 	 �      3    , "p  �� .(  �� .(  ި "p  ި "p  ��      3    , � � �� � �� 2� � 2� � �      3    , l� � x@ � x@ � l� � l� �      3    , ˈ � �@ � �@ )  ˈ )  ˈ �      3    , T� J `� J `� m4 T� m4 T� J      3    , v� �� �H �� �H ø v� ø v� ��      3    , @ 	u� � 	u� � 
k� @ 
k� @ 	u�      3    , X� 
`@ dH 
`@ dH � X� � X� 
`@      3    , �t �� �, �� �, �� �t �� �t ��      3    , k� �� wd �� wd �� k� �� k� ��      3    , *�  �0 *��  �0 *�� H  *� H  *�  �0      3    , `� [| l` [| l` "� `� "� `� [|      3    , �� 
�x �d 
�x �d � �� � �� 
�x      3    , $l  �� $$  �� $$  ި $l  ި $l  ��      3    , v� �4 �� �4 �� �� v� �� v� �4      3    , , ��  � ��  � �� , �� , ��      3    , '�� %�� '�@ %�� '�@ &� '�� &� '�� %��      3    , P $�� " $�� " %�t P %�t P $��      3    , �P �< � �< � !� �P !� �P �<      3    , 
�| t 
�4 t 
�4 6� 
�| 6� 
�| t      3    , � !�� �� !�� �� " � " � !��      3    , �| !�� �4 !�� �4 " �| " �| !��      3    , �t �| �, �| �, �4 �t �4 �t �|   	   3    !    �  &=  � &=  ��      3    , 'b 	� 'm� 	� 'm� :L 'b :L 'b 	�      3    , 'ǘ �� '�P �� '�P a 'ǘ a 'ǘ ��      3    , d� �4 p� �4 p� 	bX d� 	bX d� �4      3    , �� �4 �� �4 �� 	bX �� 	bX �� �4      3    ,    	�x  � 	�x  � ��    ��    	�x      3    , &5@ t� &@� t� &@� �� &5@ �� &5@ t�      3    , &�l �� '
$ �� '
$ 0  &�l 0  &�l ��      3    , 	�� � 	�` � 	�` 2� 	�� 2� 	�� �      3    ,  �� ��  Ơ ��  Ơ �0  �� �0  �� ��      3    , !,  �0 !�  �0 !� �� !, �� !,  �0      3    , 
h i� 
s� i� 
s� � 
h � 
h i�      3    , '� C� '�l C� '�l vp '� vp '� C�      3    , ,k �4 ,v� �4 ,v� �� ,k �� ,k �4      3    , �  v� θ v� θ @( �  @( �  v�      3    , �� $ ܈ $ ܈ :L �� :L �� $      3    , #l �� /$ �� /$ ø #l ø #l ��      3    , �� \ ݨ \ ݨ 6� �� 6� �� \      3    , �� \ �� \ �� 6� �� 6� �� \      3    , ̀ %�$ �8 %�$ �8 %�t ̀ %�t ̀ %�$      3    , � !� $d !� $d !�d � !�d � !�      3    , '�0 	bX '�� 	bX '�� 	� '�0 	� '�0 	bX      3    , %=4  �0 %H�  �0 %H� ! %=4 ! %=4  �0      3    , *6�  �x *B\  �x *B\ X *6� X *6�  �x      3    , 	�� !�, 	�P !�, 	�P !�d 	�� !�d 	�� !�,      3    , +�X !�< +� !�< +� !�d +�X !�d +�X !�<      3    , ,�� !�< ,�h !�< ,�h !�d ,�� !�d ,�� !�<      3    , 
90 %�� 
D� %�� 
D� &$ 
90 &$ 
90 %��      3    , 	�P %�� 	� %�� 	� &$ 	�P &$ 	�P %��      3    , 
��  �0 
�H  �0 
�H �� 
�� �� 
��  �0      3    ,  4$ t�  ?� t�  ?� �  4$ �  4$ t�      3    , 9� �, Ex �, Ex �T 9� �T 9� �,      3    , �$ �d �� �d �� �  �$ �  �$ �d      3    , ٜ !�< �T !�< �T !�d ٜ !�d ٜ !�<      3    , �4 a| �� a| �� !� �4 !� �4 a|      3    , D \ O� \ O� 6� D 6� D \      3    , "l �� "($ �� "($ �4 "l �4 "l ��      3    , %�d � %� � %� �� %�d �� %�d �      3    , �4  �0 ��  �0 �� 8� �4 8� �4  �0      3    , ��  �   �  8� �� 8� ��  �      3    , 0�  �0 <d  �0 <d �� 0� �� 0�  �0      3    , m8 �( x� �( x� �� m8 �� m8 �(      3    , �� �� �l �� �l �\ �� �\ �� ��      3    , �t K0 �, K0 �, nX �t nX �t K0      3    , �l � �$ � �$ L$ �l L$ �l �      3    , %�� � %׀ � %׀ 7� %�� 7� %�� �      3    , � |� )h |� )h �� � �� � |�      3    , X |�  |�  �� X �� X |�      3    , �$  �x ��  �x �� 6  �$ 6  �$  �x      3    , "5� \ "A� \ "A� 6� "5� 6� "5� \      3    , "?� `< "KL `< "KL  "?�  "?� `<   	   3    !    �  (c� I� (c� Ml      3    , 	J� i� 	V� i� 	V� � 	J� � 	J� i�      3    , !&T $ !2 $ !2 F !&T F !&T $      3    , )P, 	u� )[� 	u� )[� 	� )P, 	� )P, 	u�      3    , �| �� 4 �� 4 ø �| ø �| ��      3    , op �� {( �� {( ø op ø op ��      3    , 80 %�L C� %�L C� %�P 80 %�P 80 %�L      3    , $հ 	u� $�h 	u� $�h �� $հ �� $հ 	u�      3    , %T� �( %`\ �( %`\ �P %T� �P %T� �(      3    , � %$ �� %$ �� %�, � %�, � %$      3    , �d C� � C� � �  �d �  �d C�      3    , \x 	� h0 	� h0 6  \x 6  \x 	�      3    , ,*� �� ,6\ �� ,6\ �� ,*� �� ,*� ��      3    , +�� �D +�� �D +�� �l +�� �l +�� �D      3    , � �� �P �� �P ø � ø � ��      3    , 
�| �� 
�4 �� 
�4 ø 
�| ø 
�| ��      3    , %� o, %T o, %T @( %� @( %� o,      3    , "�  $ #� $ #� :L "�  :L "�  $      3    , $� t� $�x t� $�x �� $� �� $� t�      3    , �0 %�� �� %�� �� &$ �0 &$ �0 %��      3    , ʬ � �d � �d 0  ʬ 0  ʬ �      3    ,  !�< � !�< � !�d  !�d  !�<      3    , �� !�� �� !�� �� "�� �� "�� �� !��      3    , �| �d �4 �d �4 �� �| �� �| �d      3    , !� t� !�� t� !�� �x !� �x !� t�      3    , �p  �� �(  �� �(  ި �p  ި �p  ��      3    , ��  �X �@  �X �@  �H ��  �H ��  �X      3    , !b�  �� !n�  �� !n�  ި !b�  ި !b�  ��      3    , ![  �0 !f�  �0 !f� �� ![ �� ![  �0      3    , 	�< |� 	�� |� 	�� �� 	�< �� 	�< |�      3    , � |� �\ |� �\ �� � �� � |�      3    , H< �, S� �, S� �T H< �T H< �,      3    , �0 �, �� �, �� �T �0 �T �0 �,      3    , �� !, �8 !, �8 m4 �� m4 �� !,      3    , �X J � J � m4 �X m4 �X J      3    ,  �  !��  ¸ !��  ¸ "��  �  "��  �  !��      3    , &�0 t� &�� t� &�� �� &�0 �� &�0 t�      3    , U� �d a8 �d a8 ( U� ( U� �d      3    , μ L �t L �t �� μ �� μ L      3    , ,�` %�� ,� %�� ,� &$ ,�` &$ ,�` %��      3    , �� i� ݬ i� ݬ � �� � �� i�      3    , � !�< � !�< � !�d � !�d � !�<      3    , � !�� !t !�� !t "$< � "$< � !��      3    , )JP  �� )V  �� )V  ި )JP  ި )JP  ��      3    , )R   �0 )]�  �0 )]� �p )R  �p )R   �0      3    ,   �P  � �P  � <d   <d   �P      3    , � �� �H �� �H �� � �� � ��      3    , ~� �< �� �< ��  ~�  ~� �<      3    , � �� �� �� ��  �  � ��      3    , O� �� [8 �� [8 m� O� m� O� ��      3    , 	�  � 	�� � 	�� �� 	�  �� 	�  �      3    , :p #�t F( #�t F( $� :p $� :p #�t      3    , +�  �4 +�� �4 +�� �� +�  �� +�  �4      3    , +D, �� +O� �� +O� a +D, a +D, ��      3    , +� i� 7� i� 7� � +� � +� i�      3    ,  G� 	u�  Sd 	u�  Sd 
�H  G� 
�H  G� 	u�      3    , #�H !8 #�  !8 #�  !�d #�H !�d #�H !8      3    , "�� #�� "�� #�� "�� #�� "�� #�� "�� #��      3    , 	`d �L 	l �L 	l :L 	`d :L 	`d �L      3    , ;l �L G$ �L G$ :L ;l :L ;l �L      3    , -A� �� -M� �� -M� �� -A� �� -A� ��      3    , -e �, -p� �, -p� Ӝ -e Ӝ -e �,      3    , �< �d �� �d �� �� �< �� �< �d      3    ,  �� �d  � �d  � ��  �� ��  �� �d      3    , ( �  3� �  3� �P ( �P ( �       3    , z 
A  �� 
A  �� �� z �� z 
A       3    , �, ?x �� ?x �� C< �, C< �, ?x      3    , 'w�  �0 '�<  �0 '�< � 'w� � 'w�  �0      3    , 
p $�� ( $�� ( %�t 
p %�t 
p $��      3    , �� #�t �@ #�t �@ $� �� $� �� #�t      3    , &1X � &= � &= <d &1X <d &1X �      3    , .L �� : �� : '0 .L '0 .L ��      3    , )�� �� )�X �� )�X �P )�� �P )�� ��      3    , �4 � �� � �� )  �4 )  �4 �      3    , {p  �� �(  �� �(  ި {p  ި {p  ��      3    , � 	u� � 	u� � Rp � Rp � 	u�      3    , , F� � F� � :L , :L , F�      3    , - �� -� �� -� �d - �d - ��      3    , �  M� ڸ M� ڸ �\ �  �\ �  M�      3    , �| ̤ �4 ̤ �4 a �| a �| ̤      3    , "�D � "�� � "�� /D "�D /D "�D �      3    , &| �| 24 �| 24 �� &| �� &| �|      3    , �  �| �� �| �� �� �  �� �  �|      3    , � 	u� @ 	u� @ 
k� � 
k� � 	u�      3    , 7� M� C� M� C� p� 7� p� 7� M�      3    , �| ?x �4 ?x �4 �� �| �� �| ?x      3    , 
D� �� 
P� �� 
P� #  
D� #  
D� ��      3    , (�� |� (�� |� (�� �� (�� �� (�� |�      3    , ( < |� (� |� (� �� ( < �� ( < |�      3    , � �� d �� d � � � � ��      3    , �� �� �� �� �� @ �� @ �� ��      3    , #nP � #z � #z �� #nP �� #nP �      3    , � L �� L �� {L � {L � L      3    , p� 4P |l 4P |l 0  p� 0  p� 4P      3    , `� � l� � l� �0 `� �0 `� �      3    , �h ET �  ET �  �� �h �� �h ET      3    , ,� �( 8x �( 8x �P ,� �P ,� �(      3    ,  �� $פ  �l $פ  �l %�t  �� %�t  �� $פ      3    , �� � �P � �P 2� �� 2� �� �      3    , '�l �� ($ �� ($ u� '�l u� '�l ��      3    , '�� �d '� �d '� K, '�� K, '�� �d      3    , � #�� �h #�� �h #�� � #�� � #��      3    , 0� #�� <� #�� <� #�� 0� #�� 0� #��      3    , �� M� �� M� �� l �� l �� M�      3    , e� � qh � qh a e� a e� �      3    , z� ֌ �x ֌ �x a z� a z� ֌      3    , 0� � <d � <d �� 0� �� 0� �      3    , �� 	?0 ˨ 	?0 ˨ 	bX �� 	bX �� 	?0      3    , up Z� �( Z� �( 	bX up 	bX up Z�      3    , � S� d S� d :L � :L � S�      3    , Q, � \� � \� _� Q, _� Q, �      3    , �� 	� ۔ 	� ۔ � �� � �� 	�      3    , �d `< � `< � �l �d �l �d `<      3    , !�h `< !�  `< !�   !�h  !�h `<      3    , o� �� {P �� {P �� o� �� o� ��      3    , �� �� �` �� �` �� �� �� �� ��      3    , �| �l �4 �l �4 a �| a �| �l      3    , ڼ 7� �t 7� �t �p ڼ �p ڼ 7�      3    , a� � m8 � m8 �4 a� �4 a� �      3    , ]� � it � it �4 ]� �4 ]� �      3    , x K0 �� K0 �� �� x �� x K0      3    , '� i� '#� i� '#� �� '� �� '� i�      3    , )� �� )�H �� )�H ø )� ø )� ��      3    , � � � � � 7� � 7� � �      3    , 1� �x =` �x =` 7� 1� 7� 1� �x      3    , �l �� �$ �� �$ �� �l �� �l ��      3    , �� �� �� �� �� ̨ �� ̨ �� ��      3    , ~� �� �< �� �< 5� ~� 5� ~� ��      3    , " 
�h -� 
�h -� �� " �� " 
�h      3    , �� 	u� �@ 	u� �@ 
�  �� 
�  �� 	u�      3    , "�� %�L "� %�L "� %�t "�� %�t "�� %�L      3    , !�  %�L !�� %�L !�� %�t !�  %�t !�  %�L      3    , �� Z� �� Z� �� 	n �� 	n �� Z�   	   3    !    �  2� Q 2� T�      3    , ,�� C� ,Ԑ C� ,Ԑ �0 ,�� �0 ,�� C�      3    , ,g0 �� ,r� �� ,r� ø ,g0 ø ,g0 ��      3    ,   �d � �d � t   t   �d      3    , r� hT ~� hT ~� �� r� �� r� hT      3    , +&� �� +2� �� +2� �0 +&� �0 +&� ��      3    , ''p o, '3( o, '3( :L ''p :L ''p o,      3    , �< �< �� �< �� !0 �< !0 �< �<      3    , q@ �( |� �( |� �P q@ �P q@ �(      3    , �, |� �� |� �� �� �, �� �, |�      3    ,  �� J  �� J  �� g4  �� g4  �� J      3    , �l "b� �$ "b� �$ #�� �l #�� �l "b�      3    , � , �� , �� �� � �� � ,      3    , 	�4 C� 	�� C� 	�� `� 	�4 `� 	�4 C�      3    , �� U �L U �L 
� �� 
� �� U      3    , �� �� �x �� �x 	bX �� 	bX �� ��      3    , � ?x �t ?x �t �x � �x � ?x      3    , 
� v� 
�� v� 
�� :L 
� :L 
� v�      3    ,  � � � � )   )   �      3    , �| � �4 � �4 �0 �| �0 �| �      3    , � �  t �  t �� � �� � �       3    , �4 � �� � �� �0 �4 �0 �4 �      3    , �H � �  � �  �0 �H �0 �H �      3    , �� =� 8 =� 8 a �� a �� =�      3    , �� �d �� �d �� �� �� �� �� �d      3    , -Q�  � -]H  � -]H !�d -Q� !�d -Q�  �      3    , *�\ � *� � *�  *�\  *�\ �      3    ,  h J   J   �l  h �l  h J      3    , P �<  �<  !� P !� P �<      3    , �X K0 � K0 � nX �X nX �X K0      3    , 5� =� AH =� AH a 5� a 5� =�      3    , nX =� z =� z a nX a nX =�      3    , l� #�t x� #�t x� $� l� $� l� #�t      3    , ,� �� 8x �� 8x � ,� � ,� ��      3    , $`� � $l8 � $l8 �� $`� �� $`� �      3    , ,4 � ,� � ,� < ,4 < ,4 �      3    , -� $ -$� $ -$� :L -� :L -� $      3    , %q� ȼ %}� ȼ %}� a %q� a %q� ȼ      3    , �� �| ̄ �| ̄ �� �� �� �� �|      3    , Ĵ �, �l �, �l �T Ĵ �T Ĵ �,      3    , �T %o� � %o� � %�t �T %�t �T %o�      3    , %< � 0� � 0� I� %< I� %< �      3    , M� � Yh � Yh )  M� )  M� �      3    , #� �� /H �� /H N@ #� N@ #� ��      3    , 
T� K0 
`@ K0 
`@ �t 
T� �t 
T� K0      3    ,  � *� � *� 	bX  	bX  �      3    , 	q� i� 	}� i� 	}� � 	q� � 	q� i�      3    , W� 	?0 cL 	?0 cL 	bX W� 	bX W� 	?0      3    , :$ 	u� E� 	u� E� 
�p :$ 
�p :$ 	u�      3    , �� �  �8 �  �8 �P �� �P �� �       3    , � d� �� d� �� �� � �� � d�      3    , �� �� �� �� �� u� �� u� �� ��      3    , "tP i� "� i� "� �4 "tP �4 "tP i�      3    , !� t� !� t� !� �� !� �� !� t�      3    , )0� �� )<� �� )<� �� )0� �� )0� ��      3    , �� � �T � �T ,� �� ,� �� �      3    , �� �d �T �d �T �4 �� �4 �� �d      3    , (N\  �0 (Z  �0 (Z H  (N\ H  (N\  �0      3    ,  r� � r� � 0   0   r�      3    ,  r� � r� � 0   0   r�      3    , S  �, ^� �, ^� +� S  +� S  �,      3    , )� d� 5� d� 5� �� )� �� )� d�      3    , �� M� �x M� �x p� �� p� �� M�      3    , � � �� � �� �� � �� � �      3    , � �t $� �t $� �T � �T � �t      3    , %�p M� %�( M� %�( j� %�p j� %�p M�      3    , � %�L �d %�L �d %�t � %�t � %�L      3    , �� %�L � %�L � %�t �� %�t �� %�L      3    , *�@ t� *�� t� *�� � *�@ � *�@ t�      3    , � � *� � *� 2� � 2� � �      3    , C� 0� O� 0� O� 6� C� 6� C� 0�      3    , 4 4P � 4P � 0  4 0  4 4P      3    , �, �� �� �� �� � �, � �, ��      3    , � �� �� �� �� � � � � ��      3    , Y$ i� d� i� d� � Y$ � Y$ i�      3    , =� i� I� i� I� � =� � =� i�      3    , )JP �d )V �d )V � )JP � )JP �d      3    , &  �� &!� �� &!� � &  � &  ��      3    , 	N� #�t 	Z� #�t 	Z� $� 	N� $� 	N� #�t      3    , �d $ � � $ � � %�P �d %�P �d $ �      3    , 
�< �< 
�� �< 
�� !�� 
�< !�� 
�< �<      3    , �4 �� �� �� �� �� �4 �� �4 ��      3    ,  �< t�  �� t�  �� ��  �< ��  �< t�      3    ,  zt ��  �, ��  �, }   zt }   zt ��      3    ,  t� 
ш  �P 
ш  �P �  t� �  t� 
ш      3    , %;@ 	?0 %F� 	?0 %F� 	bX %;@ 	bX %;@ 	?0      3    , � ~@ �� ~@ �� 7� � 7� � ~@      3    , �|  �� �4  �� �4  ި �|  ި �|  ��      3    , �0 O� �� O� �� �0 �0 �0 �0 O�      3    , �l  �0 �$  �0 �$ �� �l �� �l  �0      3    ,  � 	u� ,X 	u� ,X 
�  � 
�  � 	u�      3    , U8 	�� `� 	�� `� � U8 � U8 	��      3    , pL K0 | K0 | 
%� pL 
%� pL K0      3    , �| 
� �4 
� �4 � �| � �| 
�      3    , �< t� �� t� �� �P �< �P �< t�      3    , !  !�L  !�L �T ! �T !       3    , � �, �L �, �L �$ � �$ � �,      3    , �� 6� �� 6� �� 6� �� 6� �� 6�      3    , �� !�< �� !�< �� !�d �� !�d �� !�<      3    , �� %�� � %�� � &$ �� &$ �� %��      3    , �@ %�� �� %�� �� &$ �@ &$ �@ %��      3    , ɐ J �H J �H m4 ɐ m4 ɐ J      3    , Y� �4 e� �4 e� B< Y� B< Y� �4      3    , .X �� . �� . ø .X ø .X ��      3    , *@ � *(� � *(� �0 *@ �0 *@ �      3    , oP !�� { !�� { " oP " oP !��      3    , ֐  � �H  � �H �l ֐ �l ֐  �      3    , �P �, � �, � �T �P �T �P �,      3    , 
� �D 
8 �D 
8 �l 
� �l 
� �D      3    , ,$� M� ,0� M� ,0� j� ,$� j� ,$� M�      3    , -�| L� .4 L� .4 6� -�| 6� -�| L�      3    , *0� x *<� x *<� �P *0� �P *0� x      3    , .� S� :l S� :l :L .� :L .� S�      3    , )�l t� )�$ t� )�$ �� )�l �� )�l t�      3    , )�� �| )�� �| )�� �� )�� �� )�� �|      3    , &f  � &q�  � &q� !�@ &f !�@ &f  �      3    , #`� "�D #l\ "�D #l\ #�� #`� #�� #`� "�D      3    , *� �< 6� �< 6� �d *� �d *� �<      3    , !zP 	� !� 	� !� B< !zP B< !zP 	�      3    , �0 %�� �� %�� �� &3L �0 &3L �0 %��      3    , �H %�� �  %�� �  &3L �H &3L �H %��      3    , e� 	 q� 	 q� 	bX e� 	bX e� 	      3    , e� 	 q@ 	 q@ 	bX e� 	bX e� 	      3    , e� !�� q� !�� q� "Gd e� "Gd e� !��      3    , e� !`� q� !`� q� !�d e� !�d e� !`�      3    , )� �� )#@ �� )#@ � )� � )� ��      3    , )� � *� � *� �0 )� �0 )� �      3    ,  a !�<  l� !�<  l� !�d  a !�d  a !�<      3    , ~<  �� ��  �� ��  ި ~<  ި ~<  ��      3    , 7� 	u� C� 	u� C� 	� 7� 	� 7� 	u�      3    , L� 	�` XH 	�` XH � L� � L� 	�`      3    , X $   $   :L X :L X $      3    , ې $ �H $ �H :L ې :L ې $      3    , � 	?0 � 	?0 � 	bX � 	bX � 	?0      3    , !, 	?0 ,� 	?0 ,� 	bX !, 	bX !, 	?0      3    , � � d � d �P � �P � �      3    , AD 	u� L� 	u� L� 
�0 AD 
�0 AD 	u�      3    , +M� 	u� +Y� 	u� +Y� 	� +M� 	� +M� 	u�      3    , )� 	j( )�H 	j( )�H 	� )� 	� )� 	j(      3    , !� t� -t t� -t G� !� G� !� t�      3    , �� ;� �� ;� �� �� �� �� �� ;�      3    , �� J �� J �� g4 �� g4 �� J      3    , � � �l � �l 6� � 6� � �      3    , v� K0 �� K0 �� fd v� fd v� K0      3    , �l ?x �$ ?x �$ �� �l �� �l ?x      3    , � \ �� \ �� 	bX � 	bX � \      3    , l �� $ �� $ �X l �X l ��      3    , �p � �( � �( 0  �p 0  �p �      3    , �  �0 *d  �0 *d �� � �� �  �0      3    , � >� ` >� ` �P � �P � >�      3    , N� F� Z` F� Z` � N� � N� F�      3    , �( 
�� �� 
�� �� � �( � �( 
��      3    , "l 	u� "($ 	u� "($ 	� "l 	� "l 	u�      3    , !� �8 -� �8 -� 7� !� 7� !� �8      3    , W, C� b� C� b� �  W, �  W, C�      3    , �l  u0 �$  u0 �$  ި �l  ި �l  u0      3    , ��  �X ��  �X ��  ި ��  ި ��  �X      3    , �(  �X ��  �X ��  ި �(  ި �(  �X      3    , )�� %�t )�X %�t )�X &$ )�� &$ )�� %�t      3    , �P d� � d� � �� �P �� �P d�      3    , �� d� � d� � �� �� �� �� d�      3    , *��  �0 *ޜ  �0 *ޜ �� *�� �� *��  �0      3    , *�� �� *�8 �� *�8 � *�� � *�� ��      3    , 9,  �0 D�  �0 D� �� 9, �� 9,  �0      3    , f  �� q�  �� q�  ި f  ި f  ��      3    , �� �� � �� � 	bX �� 	bX �� ��      3    , " 	u� -� 	u� -� 	�0 " 	�0 " 	u�      3    , �� 	u� �� 	u� �� 	�0 �� 	�0 �� 	u�      3    , � � t � t 7� � 7� � �      3    , I� � U� � U� L( I� L( I� �      3    , N@ � Y� � Y� L( N@ L( N@ �      3    , �| ;l �4 ;l �4 	bX �| 	bX �| ;l      3    , �, K0 �� K0 �� G$ �, G$ �, K0      3    , ϴ #�t �l #�t �l $�� ϴ $�� ϴ #�t      3    , $=X #�� $I #�� $I #�� $=X #�� $=X #��      3    , Ҥ $ �\ $ �\ :L Ҥ :L Ҥ $      3    , �� $ �d $ �d :L �� :L �� $      3    , PT � \ � \ I� PT I� PT �      3    , ,�H � ,�  � ,�  2� ,�H 2� ,�H �      3    , +�` � +� � +� 2� +�` 2� +�` �      3    , t� � �T � �T  t�  t� �      3    , f� �� r` �� r` 4 f� 4 f� ��      3    , &�P t� &� t� &� �$ &�P �$ &�P t�      3    , (� i� (�l i� (�l 6� (� 6� (� i�      3    ,  � !�  � !�  � !�@  � !�@  � !�      3    , %�� �� &l �� &l m� %�� m� %�� ��      3    , !� �P !"l �P !"l �l !� �l !� �P      3    , -:  #�t -E� #�t -E� $� -:  $� -:  #�t      3    , ̀ !�< �8 !�< �8 !�d ̀ !�d ̀ !�<      3    , Q, !�< \� !�< \� !�d Q, !�d Q, !�<      3    , U� 	� a� 	� a� _� U� _� U� 	�      3    , $�0 K0 $�� K0 $�� �� $�0 �� $�0 K0      3    , �� 
�P �� 
�P �� �� �� �� �� 
�P      3    , �� 	Ӡ �� 	Ӡ �� 
� �� 
� �� 	Ӡ      3    , �� 	u� 	� 	u� 	� 
o� �� 
o� �� 	u�      3    , y� K0 �� K0 �� �� y� �� y� K0      3    , +�H C� +�  C� +�  f� +�H f� +�H C�      3    , +�H _  +�  _  +�  �X +�H �X +�H _       3    , '�( 
� '�� 
� '�� C` '�( C` '�( 
�      3    , -�, � -�� � -�� 7� -�, 7� -�, �      3    , �� 	?0 �| 	?0 �| 	bX �� 	bX �� 	?0      3    , �8 
= �� 
= �� � �8 � �8 
=      3    , � %�D 't %�D 't &$ � &$ � %�D      3    , �� eD �� eD �� l� �� l� �� eD      3    , (%X 	� (1 	� (1 :L (%X :L (%X 	�      3    , (%X M� (1 M� (1 �L (%X �L (%X M�      3    , (�< �� )� �� )�  (�<  (�< ��      3    , ,�� |� ,�� |� ,�� �� ,�� �� ,�� |�      3    , ,�� �< ,�t �< ,�t  � ,��  � ,�� �<      3    , )6� !�� )B� !�� )B� " )6� " )6� !��      3    , �� d� ˨ d� ˨ �� �� �� �� d�      3    , �� d� �P d� �P �� �� �� �� d�      3    , �� �� �� �� ��  ��  �� ��      3    , � Ӝ &� Ӝ &�  �  � Ӝ      3    , T` , ` , ` �� T` �� T` ,      3    , !b� �� !n� �� !n� '0 !b� '0 !b� ��      3    , &  	u� &!� 	u� &!� 
)� &  
)� &  	u�      3    , &�� Y� &�� Y� &�� �0 &�� �0 &�� Y�      3    , �� � �p � �p 7� �� 7� �� �      3    , �� z� � z� � j� �� j� �� z�      3    , ר �( �` �( �` 7� ר 7� ר �(      3    , Z�  �0 f`  �0 f` 8� Z� 8� Z�  �0      3    , 6� �� Bd �� Bd ø 6� ø 6� ��      3    , �� �� � �� � ̨ �� ̨ �� ��      3    , �� C� �8 C� �8 7� �� 7� �� C�      3    , )�� K0 )�@ K0 )�@ �� )�� �� )�� K0      3    , #^� � #jh � #jh )  #^� )  #^� �      3    , )�� � )�X � )�X _� )�� _� )�� �      3    , (� B� 4l B� 4l �P (� �P (� B�      3    , M� �, Yd �, Yd �D M� �D M� �,      3    ,  �l b�  �$ b�  �$ hX  �l hX  �l b�      3    , #�@ �� #�� �� #�� ̨ #�@ ̨ #�@ ��      3    , �` �4 � �4 � �� �` �� �` �4      3    , � J �� J �� m4 � m4 � J      3    , &�� �� &�� �� &�� 6� &�� 6� &�� ��      3    , &i� � &u� � &u� � &i� � &i� �      3    , 
�L 1 
� 1 
� �P 
�L �P 
�L 1      3    , =� � I� � I� oP =� oP =� �      3    , Ș i� �P i� �P � Ș � Ș i�      3    , ��  �0 ��  �0 �� 8� �� 8� ��  �0      3    , $`� �, $l8 �, $l8 k� $`� k� $`� �,      3    , '>� � 'J� � 'J� �� '>� �� '>� �      3    , )uH K0 )�  K0 )�  	G  )uH 	G  )uH K0      3    , �` C� � C� � �� �` �� �` C�      3    , 	�� |( 	�� |( 	�� 7� 	�� 7� 	�� |(      3    , 
�� 	?0 8 	?0 8 	bX 
�� 	bX 
�� 	?0      3    , � K0 �� K0 �� hX � hX � K0      3    , �0 K0 � K0 � nX �0 nX �0 K0      3    , $�P =� $� =� $� a $�P a $�P =�      3    , %5d �� %A �� %A � %5d � %5d ��      3    , "/� ?x ";� ?x ";� �� "/� �� "/� ?x      3    , !�P � " � " 	bX !�P 	bX !�P �      3    , � � t � t 7� � 7� � �      3    , ֈ � �@ � �@ 7� ֈ 7� ֈ �      3    , �p t� 
( t� 
( �� �p �� �p t�      3    , m� G� y| G� y| C� m� C� m� G�      3    , &�� �\ 'H �\ 'H �� &�� �� &�� �\      3    , (�� � (�� � (�� �4 (�� �4 (�� �      3    , �P C� � C� � f� �P f� �P C�      3    , �P �� � �� � � �P � �P ��      3    , !`� |� !l� |� !l� �� !`� �� !`� |�      3    , � |� �� |� �� �� � �� � |�      3    , -I� �� -Ux �� -Ux �� -I� �� -I� ��      3    , " =� "� =� "� a " a " =�      3    , $� !�< $�� !�< $�� !�d $� !�d $� !�<      3    , 
1` K0 
= K0 
= 	'� 
1` 	'� 
1` K0      3    , �d � � � � � �d � �d �      3    , � d� �� d� �� �� � �� � d�      3    , � �h �� �h �� 7� � 7� � �h      3    , �T �� � �� � �� �T �� �T ��      3    , �� 	u� �H 	u� �H 	� �� 	� �� 	u�      3    , �$ � �� � �� �4 �$ �4 �$ �      3    , C� �� O� �� O�  C�  C� ��      3    , �H � �  � �  F$ �H F$ �H �      3    , �H �T �  �T �  �4 �H �4 �H �T      3    , xd \� � \� � 	A$ xd 	A$ xd \�      3    , %< J 0� J 0� g4 %< g4 %< J      3    , 4P �4 @ �4 @ �� 4P �� 4P �4      3    ,  � #ټ  �t #ټ  �t $+�  � $+�  � #ټ      3    , !;� #�� !G� #�� !G� #�� !;� #�� !;� #��      3    , *�� �� *ڴ �� *ڴ  *��  *�� ��      3    , +� �� +�� �� +��  +�  +� ��      3    ,  D �< � �< � �  D �  D �<      3    , 
 �4 � �4 � , 
 , 
 �4      3    , X� %$ d� %$ d� %�t X� %�t X� %$      3    , � #�t �� #�t �� %!� � %!� � #�t      3    , �� =� �8 =� �8 a �� a �� =�      3    , �l =� �$ =� �$ f� �l f� �l =�      3    , �( � �� � �� �� �( �� �( �      3    , �h M� �  M� �  p� �h p� �h M�      3    , *�  �� +� �� +� � *�  � *�  ��      3    , "� �( "�� �( "�� �, "� �, "� �(      3    , �  	׈ Ը 	׈ Ը � �  � �  	׈      3    , P J [� J [� m4 P m4 P J      3    , � J � J � m4 � m4 � J      3    , h J   J   m4 h m4 h J      3    , 'P �D 3 �D 3 �l 'P �l 'P �D      3    , >0 �� I� �� I� /D >0 /D >0 ��      3    , $"  �� $-� �� $-� �� $"  �� $"  ��      3    , !�H M� !�  M� !�  �� !�H �� !�H M�      3    , �� #�� � #�� � #�� �� #�� �� #��      3    , ϐ #�� �H #�� �H #�� ϐ #�� ϐ #��      3    , �� + �8 + �8 6� �� 6� �� +      3    , �  �� �t  �� �t #�� � #�� �  ��      3    , 	�� "� 	�� "� 	�� #� 	�� #� 	�� "�      3    , U� %�$ a� %�$ a� %� U� %� U� %�$      3    , !�� �� !�� �� !�� �� !�� �� !�� ��      3    ,  �� ��  �� ��  �� ��  �� ��  �� ��      3    , *� � *| � *| �� *� �� *� �      3    , **� J *6� J *6� �� **� �� **� J      3    , {P �� � �� � 5� {P 5� {P ��      3    , 
V|  �x 
b4  �x 
b4 <h 
V| <h 
V|  �x      3    ,  �P \ !	 \ !	 	bX  �P 	bX  �P \      3    , &P� i� &\P i� &\P � &P� � &P� i�      3    , 	j( �, 	u� �, 	u� +� 	j( +� 	j( �,      3    , �� �D 	
t �D 	
t �l �� �l �� �D      3    , "�p #�� "�( #�� "�( #�� "�p #�� "�p #��      3    , %�H #�t %�  #�t %�  $+� %�H $+� %�H #�t      3    , "�� $C4 "�X $C4 "�X %�, "�� %�, "�� $C4      3    , �| $�� 4 $�� 4 %�P �| %�P �| $��      3    , �, �D �� �D �� �l �, �l �, �D      3    , �P �d � �d � w� �P w� �P �d      3    , eh J q  J q  m4 eh m4 eh J      3    , 1� �< =� �< =� 4 1� 4 1� �<      3    , # 0 � #+� � #+� )  # 0 )  # 0 �      3    , , 84  � 84  � l� , l� , 84      3    , �P  �0 �  �0 � X �P X �P  �0      3    , Z�  �� f�  �� f�  ި Z�  ި Z�  ��      3    , S� C� _D C� _D �p S� �p S� C�      3    , Z� ^� fd ^� fd 	�0 Z� 	�0 Z� ^�      3    , $l � $$ � $$ �0 $l �0 $l �      3    , '�l � ($ � ($ 7� '�l 7� '�l �      3    , (�p ;� (�( ;� (�( �� (�p �� (�p ;�      3    , �p � �( � �( �� �p �� �p �      3    , 
�� �, 8 �, 8 q� 
�� q� 
�� �,      3    , �l �� �$ �� �$ 	bX �l 	bX �l ��      3    , YH �l e  �l e  �� YH �� YH �l      3    , � B � B � � � � � B      3    , 
� =� 
�� =� 
�� f� 
� f� 
� =�      3    , i0 |� t� |� t� �� i0 �� i0 |�      3    , l� S� x` S� x` :L l� :L l� S�      3    , a T@ l� T@ l� �P a �P a T@      3    , �D Yd �� Yd �� �� �D �� �D Yd      3    , 	bX \ 	n \ 	n 6� 	bX 6� 	bX \      3    , 
)� \ 
5H \ 
5H 6� 
)� 6� 
)� \      3    , 4� >T @H >T @H m4 4� m4 4� >T      3    , �� �( � �( � �, �� �, �� �(      3    , )  �( 4� �( 4� �P )  �P )  �(      3    , �T !�� � !�� � " �T " �T !��      3    , �, �< �� �< �� !�� �, !�� �, �<      3    , #� #l #x #l #x #�� #� #�� #� #l      3    , �t M� �, M� �, l� �t l� �t M�      3    , �� t� �� t� �� $ �� $ �� t�      3    , {, �x �� �x �� 7� {, 7� {, �x      3    , 	�p � 	�( � 	�( )  	�p )  	�p �      3    , �( �\ �� �\ �� �� �( �� �( �\      3    , 	� �� 	+� �� 	+� � 	� � 	� ��      3    ,  � t� ,8 t� ,8 ��  � ��  � t�      3    , �� �� �d �� �d a �� a �� ��      3    , 	ϸ �� 	�p �� 	�p 	bX 	ϸ 	bX 	ϸ ��      3    , �< 
ɸ � 
ɸ � � �< � �< 
ɸ      3    , � �� | �� | �� � �� � ��      3    , � i, � i, � a � a � i,      3    , 
5H 4( 
A  4( 
A  a 
5H a 
5H 4(      3    , 	�� =� 	�8 =� 	�8 a 	�� a 	�� =�      3    , �H �� �  �� �  �P �H �P �H ��      3    , �� �� �� �� �� �� �� �� �� ��      3    , Rp  �0 ^(  �0 ^( X Rp X Rp  �0      3    , +| K0 +4 K0 +4 �� +| �� +| K0      3    , +| 28 +4 28 +4 7� +| 7� +| 28      3    , ��  �0 ��  �0 �� �X �� �X ��  �0      3    , ��  �0 �t  �0 �t �� �� �� ��  �0      3    , O< K0 Z� K0 Z�   O<   O< K0      3    , SH K0 _  K0 _  nX SH nX SH K0      3    , 5� !�� AD !�� AD "�� 5� "�� 5� !��      3    , 	� K0 t K0 t �� 	� �� 	� K0      3    , Y� K0 e@ K0 e@ �� Y� �� Y� K0      3    , +[� J +gT J +gT �T +[� �T +[� J      3    , +cl i� +o$ i� +o$ 6� +cl 6� +cl i�      3    , 
�� ^�  h ^�  h C< 
�� C< 
�� ^�      3    , VX e� b e� b �P VX �P VX e�      3    , � �� ` �� ` 	bX � 	bX � ��      3    , >X 	u� J 	u� J 	� >X 	� >X 	u�      3    , �� K0 �� K0 �� nX �� nX �� K0      3    , X @  @  ;� X ;� X @      3    , �� ��  d ��  d c0 �� c0 �� ��      3    , �x =� �0 =� �0 h �x h �x =�      3    , �l C� �$ C� �$ f� �l f� �l C�      3    , �� �< �� �< �� �d �� �d �� �<      3    , 	�� "�� 	�l "�� 	�l #�� 	�� #�� 	�� "��      3    , &Xh K0 &d  K0 &d  �� &Xh �� &Xh K0      3    , #�� K0 #�l K0 #�l �� #�� �� #�� K0      3    , 	X ��  ��  �� 	X �� 	X ��      3    , ]T t� i t� i �� ]T �� ]T t�      3    , &L� � &Xh � &Xh �0 &L� �0 &L� �      3    , '\, � 'g� � 'g� �0 '\, �0 '\, �      3    , #�  M� #�� M� #�� �t #�  �t #�  M�      3    , $I 	u� $T� 	u� $T� 
� $I 
� $I 	u�      3    , l� D0 x< D0 x< m4 l� m4 l� D0      3    , *�� � *�@ � *�@ V *�� V *�� �      3    , &� D0 &Ǽ D0 &Ǽ m4 &� m4 &� D0      3    , +� !�� +@ !�� +@ " +� " +� !��      3    , "�� !�� "�x !�� "�x #"$ "�� #"$ "�� !��      3    , !�  �� !"l  �� !"l !�d !� !�d !�  ��      3    , "p �| .( �| .( �4 "p �4 "p �|      3    , �` ', � ', � 6� �` 6� �` ',      3    , � M� 8 M� 8 C� � C� � M�      3    , P t� ! t� ! �� P �� P t�      3    , +<\ \ +H \ +H 6� +<\ 6� +<\ \      3    , ,W� \ ,cH \ ,cH 6� ,W� 6� ,W� \      3    ,  .H K0  :  K0  :  ��  .H ��  .H K0      3    , �� �< 	� �< 	� �� �� �� �� �<      3    , �� K0 �8 K0 �8 nX �� nX �� K0      3    , �, w  �� w  �� �0 �, �0 �, w       3    , �  �0 l  �0 l �� � �� �  �0      3    , �4 �@ �� �@ �� �0 �4 �0 �4 �@      3    , �� �� �� �� �� @ �� @ �� ��      3    , , 4P '� 4P '� 0  , 0  , 4P      3    , 'P  �� 3  �� 3  ި 'P  ި 'P  ��      3    ,   �� �  �� �  ި   ި   ��      3    , 0� Đ <` Đ <` 7� 0� 7� 0� Đ      3    , �0 �| �� �| �� �� �0 �� �0 �|      3    , �� �d �� �d �� �4 �� �4 �� �d      3    , �| |� 	4 |� 	4 �� �| �� �| |�      3    , �X |� 	 |� 	 �l �X �l �X |�      3    , #�0 \ #�� \ #�� 6� #�0 6� #�0 \      3    , � J �d J �d e � e � J      3    , '0 �� '� �� '� �4 '0 �4 '0 ��      3    , � �$ t �$ t %\ � %\ � �$      3    , �p #�� �( #�� �( $� �p $� �p #��      3    , tX � � � � �4 tX �4 tX �      3    , vp �� �( �� �( 6� vp 6� vp ��      3    , #�p � #�( � #�( �� #�p �� #�p �      3    , %�0 �8 %�� �8 %�� 0  %�0 0  %�0 �8      3    , `` �� l �� l � `` � `` ��      3    ,  �` � �` � �d  �d  �`      3    , '� �� '�H �� '�H a '� a '� ��      3    , (�$ �� )	� �� )	� a (�$ a (�$ ��      3    , $�< � $�� � $�� �4 $�< �4 $�< �      3    , &0 � &� � &� �4 &0 �4 &0 �      3    , %�� �� &` �� &` �  %�� �  %�� ��      3    , �� 	f@ �� 	f@ �� � �� � �� 	f@      3    , " C� "� C� "� �  " �  " C�      3    , �p � ( � ( 2� �p 2� �p �      3    , � %�$ �� %�$ �� %�, � %�, � %�$      3    , � �< �� �< ��  Ơ �  Ơ � �<      3    , �� %�  �8 %�  �8 &$ �� &$ �� %�       3    , D4 %�$ O� %�$ O� %�t D4 %�t D4 %�$      3    , &
H |� &  |� &  �� &
H �� &
H |�      3    , ʬ � �d � �d �4 ʬ �4 ʬ �      3    , S� � _� � _� 7� S� 7� S� �      3    ,  	�P � 	�P � ��  ��  	�P      3    , ,p� �| ,|� �| ,|� �� ,p� �� ,p� �|      3    , ,�� M� ,�8 M� ,�8 �L ,�� �L ,�� M�      3    , 5� !�� Ah !�� Ah " 5� " 5� !��      3    , -�l :l -�$ :l -�$ �l -�l �l -�l :l      3    , �l �4 �$ �4 �$ 6� �l 6� �l �4      3    , V [| a� [| a� �l V �l V [|      3    , 	?0 %o� 	J� %o� 	J� %�t 	?0 %�t 	?0 %o�      3    , $d #�t 0 #�t 0 $r $d $r $d #�t      3    , �0 "�D �� "�D �� #�� �0 #�� �0 "�D      3    , '�P � '� � '� �4 '�P �4 '�P �      3    , %�0 M� %�� M� %�� p� %�0 p� %�0 M�      3    , &� �� &#� �� &#� <` &� <` &� ��      3    , �� "� �H "� �H #�� �� #�� �� "�      3    , !�� �< !Ĉ �< !Ĉ �d !�� �d !�� �<      3    , J !�< U� !�< U� !�d J !�d J !�<      3    , �� !�< � !�< � !�d �� !�d �� !�<      3    , -�� �� -�\ �� -�\ �� -�� �� -�� ��      3    , ,�h �  ,�  �  ,�  �P ,�h �P ,�h �       3    , 3 � >� � >� �t 3 �t 3 �      3    , �� #l Ь #l Ь #�� �� #�� �� #l      3    , � � �� � �� 2� � 2� � �      3    , {P  �0 �  �0 � X {P X {P  �0      3    , �� �� �x �� �x � �� � �� ��      3    , �p  �0 (  �0 ( X �p X �p  �0   	   3    !    �P   ��  ��  �� $�� +  ,VR_LEFT_VERTICAL_BUS      3    , �H t�   t�   �� �H �� �H t�      3    , "�� �� "�p �� "�p �H "�� �H "�� ��      3    , +�� K0 +�d K0 +�d nX +�� nX +�� K0      3    , �D �� �� �� �� �4 �D �4 �D ��      3    , vp � �( � �( )  vp )  vp �      3    , �� C� �x C� �x f� �� f� �� C�      3    , S� T@ _H T@ _H �P S� �P S� T@      3    , �P � � � � )  �P )  �P �      3    , *�P �� *� �� *� �� *�P �� *�P ��      3    , !�, � !�� � !�� �� !�, �� !�, �      3    , cP %�� o %�� o &$ cP &$ cP %��      3    , ,(� � ,4h � ,4h �4 ,(� �4 ,(� �      3    , -p� M� -|� M� -|� p� -p� p� -p� M�      3    , h M�   M�   &| h &| h M�      3    , ݬ m| �d m| �d �\ ݬ �\ ݬ m|      3    , '�( �� '�� �� '�� � '�( � '�( ��      3    , '�, �� '�� �� '�� �0 '�, �0 '�, ��      3    , �� �� �| �� �| �� �� �� �� ��      3    , "� �� "� �� "� �\ "� �\ "� ��      3    , *J, �| *U� �| *U� �� *J, �� *J, �|      3    , *s0 �� *~� �� *~�  *s0  *s0 ��      3    , '�� !�< '� !�< '� !�d '�� !�d '�� !�<      3    , )�  Ĭ )|  Ĭ )| !�0 )� !�0 )�  Ĭ      3    , �$ �, �� �, �� �T �$ �T �$ �,      3    , �� ݄ �� ݄ �� �� �� �� �� ݄      3    , hX  �� t  �� t  ި hX  ި hX  ��      3    , #}�  �X #��  �X #��  ި #}�  ި #}�  �X      3    , �p �� �( �� �( �X �p �X �p ��      3    , /� , ;h , ;h !� /� !� /� ,      3    , � t� �� t� �� �� � �� � t�      3    , � �d � �d � �� � �� � �d      3    , �l 	�� �$ 	�� �$ � �l � �l 	��      3    , �4 	u� �� 	u� �� 
� �4 
� �4 	u�      3    , �X �  �  7� �X 7� �X �      3    , ., �X 9� �X 9� 7� ., 7� ., �X      3    , }   �0 ��  �0 �� X }  X }   �0      3    , w   �x ��  �x �� X w  X w   �x      3    , M� � Y� � Y� y4 M� y4 M� �      3    , "�\ !�� "� !�� "� " "�\ " "�\ !��      3    , -� J� -�� J� -�� �� -� �� -� J�      3    , .� �  .(h �  .(h �P .� �P .� �       3    , )�� � )�x � )�x �� )�� �� )�� �      3    , ,cH � ,o  � ,o  �\ ,cH �\ ,cH �      3    , �� � �� � �� 2� �� 2� �� �      3    , v� �� �� �� �� �� v� �� v� ��      3    , +4�  Ĭ +@D  Ĭ +@D !� +4� !� +4�  Ĭ      3    ,  �� !��  �� !��  �� #"$  �� #"$  �� !��      3    , �� %�� �\ %�� �\ &$ �� &$ �� %��      3    , �4 #ټ � #ټ � $R� �4 $R� �4 #ټ      3    , '< � '� � '� �� '< �� '< �      3    , $�4 |� $�� |� $�� �l $�4 �l $�4 |�      3    ,  ʈ `<  �@ `<  �@ �  ʈ �  ʈ `<      3    , "� �t .� �t .� k� "� k� "� �t      3    , E� #�� Q� #�� Q� #�� E� #�� E� #��      3    , !�� #�t !�� #�t !�� $� !�� $� !�� #�t      3    , �� eD �X eD �X p� �� p� �� eD      3    , y| \ �4 \ �4 B< y| B< y| \      3    , �@ \ � \ � 6� �@ 6� �@ \      3    , E0 !n� P� !n� P� !�d E0 !�d E0 !n�      3    , R� �, ^H �, ^H � R� � R� �,      3    , ""H ~� ".  ~� ".  :L ""H :L ""H ~�      3    , !�H x !�  x !�  �� !�H �� !�H x      3    , �� M� �� M� �� p� �� p� �� M�      3    ,  (l M�  4$ M�  4$ p�  (l p�  (l M�      3    , � � �� � �� �4 � �4 � �      3    , �  � �� � �� �4 �  �4 �  �      3    , �t � �, � �, )  �t )  �t �      3    , g� � s� � s� 2� g� 2� g� �      3    , 	Ѭ J� 	�d J� 	�d �4 	Ѭ �4 	Ѭ J�      3    , �| _D �4 _D �4 �@ �| �@ �| _D      3    , #�� 	?0 #�< 	?0 #�< 	bX #�� 	bX #�� 	?0      3    , �� �� �� �� �� �� �� �� �� ��      3    , 4� 	u� @p 	u� @p 
o� 4� 
o� 4� 	u�      3    , 4� �� @p �� @p 	bX 4� 	bX 4� ��      3    , � #�t � #�t � $� � $� � #�t      3    , m #�t x� #�t x� $� m $� m #�t      3    , -v� � -�d � -�d �l -v� �l -v� �      3    , � 	u� �D 	u� �D 
%� � 
%� � 	u�      3    , � �� �< �� �< 	bX � 	bX � ��      3    , �h  ' �   ' �   ި �h  ި �h  '      3    , p� �  |� �  |� �X p� �X p� �       3    , Y� �� e@ �� e@ #  Y� #  Y� ��      3    , S� H _@ H _@ :L S� :L S� H      3    , (� �� 4l �� 4l -0 (� -0 (� ��      3    , %�l !�< %�$ !�< %�$ !�d %�l !�d %�l !�<      3    , '�H  N  (
   N  (
   ި '�H  ި '�H  N       3    , *6� �� *B\ �� *B\ �4 *6� �4 *6� ��      3    , *>t � *J, � *J, �� *>t �� *>t �      3    , +�t �, +�, �, +�, �T +�t �T +�t �,      3    , ,d �@ , �@ , �P ,d �P ,d �@      3    , �D %�� �� %�� �� &3L �D &3L �D %��      3    , �` %�� � %�� � &3L �` &3L �` %��      3    , �, �� �� �� �� �� �, �� �, ��      3    , �� �< �� �< �� �d �� �d �� �<      3    , n4 �� y� �� y� �4 n4 �4 n4 ��      3    , fd � r � r �� fd �� fd �      3    , i0  ' t�  ' t�  ި i0  ި i0  '      3    , h�  �0 t�  �0 t� X h� X h�  �0      3    , � C� � C� � f� � f� � C�      3    , Z �� e� �� e� [< Z [< Z ��      3    , � ^� %� ^� %� ݈ � ݈ � ^�      3    , �� "� �t "� �t #�� �� #�� �� "�      3    , �@ d�  � d�  � �� �@ �� �@ d�      3    , , t� 7� t� 7� l� , l� , t�      3    , +�� \� ,� \� ,� 	bX +�� 	bX +�� \�      3    , +2� � +>P � +>P 7� +2� 7� +2� �      3    , �� %�� �t %�� �t &3L �� &3L �� %��      3    , �( � �� � �� �� �( �� �( �      3    , "Z� 
� "f� 
� "f� 7� "Z� 7� "Z� 
�      3    , $I 
� $T� 
� $T� 7� $I 7� $I 
�      3    ,  ET � ET � ��  ��  ET      3    , ", K0 -� K0 -� �� ", �� ", K0      3    , �� 	u� �\ 	u� �\ 	�8 �� 	�8 �� 	u�      3    , �� �� �P �� �P 	u� �� 	u� �� ��      3    ,  A� �,  M� �,  M� �  A� �  A� �,      3    , �` #� � #� � � �` � �` #�      3    , *c� !�< *oH !�< *oH !�d *c� !�d *c� !�<      3    , )�� !� )�� !� )�� !�@ )�� !�@ )�� !�      3    , $0 ' $%� ' $%� �T $0 �T $0 '      3    , $9p t� $E( t� $E( � $9p � $9p t�      3    , H< �� S� �� S� �� H< �� H< ��      3    , %!� �� %-� �� %-� ø %!� ø %!� ��      3    , 
7<  � 
B�  � 
B� !�@ 
7< !�@ 
7<  �      3    , FH !�� R  !�� R  "$< FH "$< FH !��      3    , 5� � A� � A� �0 5� �0 5� �      3    , K0 � V� � V� �0 K0 �0 K0 �      3    , 0� �, <� �, <� N� 0� N� 0� �,      3    , 
� C 
�� C 
�� �$ 
� �$ 
� C      3    , �l �< �$ �< �$ !� �l !� �l �<      3    , ;� %�  GH %�  GH &3L ;� &3L ;� %�       3    , �� "� �8 "� �8 #�� �� #�� �� "�      3    , =� m� I� m� I� �4 =� �4 =� m�      3    , &b, �@ &m� �@ &m� 	bX &b, 	bX &b, �@      3    , d C�  C�  �@ d �@ d C�      3    , � �� �� �� �� @ � @ � ��      3    , i0 � t� � t� 0  i0 0  i0 �      3    , d 	��  	��  � d � d 	��      3    , O� � [� � [� 	bX O� 	bX O� �      3    , 1� �� =� �� =� � 1� � 1� ��      3    , �,  �� 	�  �� 	�  �H �,  �H �,  ��      3    , 
��  �� 
�H  �� 
�H  ި 
��  ި 
��  ��      3    , 	{�  �� 	�t  �� 	�t  ި 	{�  ި 	{�  ��      3    , 
  	u� 
� 	u� 
� 
L� 
  
L� 
  	u�      3    , �� � �� � �� 7� �� 7� �� �      3    , � [| �P [| �P �� � �� � [|      3    , �d �< � �< � �d �d �d �d �<      3    , �� J �x J �x �� �� �� �� J      3    , "Ep |� "Q( |� "Q( �� "Ep �� "Ep |�      3    , #�� �< #ݤ �< #ݤ !�� #�� !�� #�� �<      3    , 	T� �� 	`d �� 	`d А 	T� А 	T� ��      3    ,  �� � �� � 0   0   ��      3    , ��  �0 �l  �0 �l X �� X ��  �0      3    , �h  �0 �   �0 �  X �h X �h  �0      3    , �< �d �� �d �� � �< � �< �d      3    , �< �D �� �D �� �� �< �� �< �D      3    , $ �D (� �D (� �l $ �l $ �D      3    , � �< �� �< �� �d � �d � �<      3    , ($ ?t (� ?t (� �$ ($ �$ ($ ?t      3    , )Y� � )e� � )e� 2� )Y� 2� )Y� �      3    , g  �� r�  �� r� !�d g !�d g  ��      3    , �X !�� � !�� � " �X " �X !��      3    , � K0 � K0 � nX � nX � K0      3    , D � )� � )� �l D �l D �      3    , �� �� �P �� �P �P �� �P �� ��      3    , � �d �8 �d �8 %� � %� � �d      3    , ��  �0 �l  �0 �l X �� X ��  �0      3    ,    �X  �  �X  �  ި    ި    �X      3    , *.� M� *:� M� *:� a *.� a *.� M�      3    , l� J x� J x� �l l� �l l� J      3    , �� �( �h �( �h �P �� �P �� �(      3    , �� �( � �( � �P �� �P �� �(      3    , & � 1� � 1� � & � & �      3    , �@   ��   �� V �@ V �@        3    , �d !�\ � !�\ � #�� �d #�� �d !�\      3    , �4 #�t �� #�t �� $+� �4 $+� �4 #�t      3    , �� �� ƨ �� ƨ �� �� �� �� ��      3    , "P � . � . 0  "P 0  "P �      3    , )�  C� )�� C� )�� � )�  � )�  C�      3    , )y0 �� )�� �� )�� 7� )y0 7� )y0 ��      3    , -> K0 -I� K0 -I� nX -> nX -> K0      3    , *�� �h *�@ �h *�@ =� *�� =� *�� �h      3    , $�� 
A  % � 
A  % � � $�� � $�� 
A       3    , �, K0 �� K0 ��   �,   �, K0      3    , &�< "^� &�� "^� &�� #�� &�< #�� &�< "^�      3    , &l !�� &$ !�� &$ "�� &l "�� &l !��      3    , $�| "�� $�4 "�� $�4 #�� $�| #�� $�| "��      3    , %� #�� %H #�� %H #�� %� #�� %� #��      3    , �� M� d M� d p� �� p� �� M�      3    , ?t M� K, M� K, p� ?t p� ?t M�      3    , Z� � fd � fd �p Z� �p Z� �      3    , �� �d �d �d �d �� �� �� �� �d      3    , g� 	� s| 	� s| V g� V g� 	�      3    , �� C� Θ C� Θ �H �� �H �� C�      3    , Nd %�L Z %�L Z %�t Nd %�t Nd %�L      3    , B� %�L N� %�L N� %�t B� %�t B� %�L      3    , � s �� s �� �0 � �0 � s      3    , |(  � ��  � ��  � |(  � |(  �      3    , W !�� b� !�� b� #�� W #�� W !��      3    , �D #�� �� #�� �� #�� �D #�� �D #��      3    , P 
�P ! 
�P ! k� P k� P 
�P      3    , "�� !�< "�@ !�< "�@ !�d "�� !�d "�� !�<      3    , +�� t� +�� t� +�� l� +�� l� +�� t�      3    , &�� �� &�d �� &�d /D &�� /D &�� ��      3    , -0 �L 8� �L 8� B< -0 B< -0 �L      3    , ��  �� �8  �� �8 !�d �� !�d ��  ��      3    , -� � 9� � 9� 5� -� 5� -� �      3    , )�H =� )�  =� )�  � )�H � )�H =�      3    , %Ә 0� %�P 0� %�P :L %Ә :L %Ә 0�      3    , -&� �� -2P �� -2P �� -&� �� -&� ��      3    , .X #� . #� . � .X � .X #�      3    , &� �@ &%� �@ &%� ;� &� ;� &� �@      3    , %� |� %�� |� %�� �0 %� �0 %� |�      3    , ,� ( ,�� ( ,�� 0  ,� 0  ,� (      3    , . �  h .,P  h .,P � . � � . �  h      3    , �� = �� = �� �l �� �l �� =      3    , "�� �d "�� �d "�� H� "�� H� "�� �d      3    , "� N@ "� N@ "� �P "� �P "� N@      3    , ,�X ȼ ,� ȼ ,� a ,�X a ,�X ȼ      3    ,  �| M�  �4 M�  �4 �L  �| �L  �| M�      3    , +@ �( +"� �( +"� �P +@ �P +@ �(      3    , 
�@ !�T 
�� !�T 
�� !�d 
�@ !�d 
�@ !�T      3    , �4 � �� � �� �� �4 �� �4 �      3    , &�P � &� � &� 0  &�P 0  &�P �      3    , &�( �� &�� �� &�� А &�( А &�( ��      3    , � �� �� �� �� ̨ � ̨ � ��      3    , &�  �� &��  �� &�� H  &� H  &�  ��      3    , |( �� �� �� ��  |(  |( ��      3    , C� L O� L O� �4 C� �4 C� L      3    , Sh ?t _  ?t _  �� Sh �� Sh ?t      3    , $d �d 0 �d 0 K, $d K, $d �d      3    , '
$ �, '� �, '� o� '
$ o� '
$ �,      3    , &{� d$ &�H d$ &�H �l &{� �l &{� d$      3    , (-( � (8� � (8� �� (-( �� (-( �      3    , )ol �� ){$ �� ){$ u� )ol u� )ol ��      3    , +�� �� +�� �� +�� /D +�� /D +�� ��      3    , +M� `< +Y� `< +Y� /D +M� /D +M� `<      3    , p� �� |� �� |� �l p� �l p� ��      3    , � � @ � @ �4 � �4 � �      3    , q  �, |� �, |� d q  d q  �,      3    , Y� C� ed C� ed �H Y� �H Y� C�      3    , (�| #ߘ (�4 #ߘ (�4 %�t (�| %�t (�| #ߘ      3    , *u$ #�t *�� #�t *�� $u� *u$ $u� *u$ #�t      3    , �� � ޤ � ޤ � �� � �� �      3    , T� �� `� �� `� �� T� �� T� ��      3    , (0 \ (� \ (� 6� (0 6� (0 \      3    , &�� \ &�� \ &�� 6� &�� 6� &�� \      3    , �  #�t ø #�t ø %�� �  %�� �  #�t      3    , #^� � #jh � #jh �0 #^� �0 #^� �      3    , �T %�L � %�L � %�t �T %�t �T %�L      3    , p( #�t {� #�t {� %� p( %� p( #�t      3    , � $ �� $ �� :L � :L � $      3    , *S� � *_� � *_� �� *S� �� *S� �      3    , �� e� �x e� �x �P �� �P �� e�      3    , �0 J �� J �� m4 �0 m4 �0 J      3    , .P J : J : m4 .P m4 .P J      3    , ]P !�D i !�D i #�� ]P #�� ]P !�D      3    , �@ $f\ �� $f\ �� %�t �@ %�t �@ $f\      3    , S� #�t _H #�t _H $�L S� $�L S� #�t      3    , � �d �� �d �� �\ � �\ � �d      3    , ,�h i� ,�  i� ,�  � ,�h � ,�h i�      3    , , i� ,$� i� ,$� � , � , i�      3    , �� Ӝ � Ӝ � �$ �� �$ �� Ӝ      3    , +�� � +ڐ � +ڐ �l +�� �l +�� �      3    , #�  �� #�� �� #�� � #�  � #�  ��      3    , "�� �� "�H �� "�H � "�� � "�� ��      3    , &  ȼ &!� ȼ &!� a &  a &  ȼ      3    ,  � f�  X f�  X ��  � ��  � f�      3    , -� � 9x � 9x � -� � -� �      3    , .S` J ._ J ._ ֬ .S` ֬ .S` J      3    , �� M� �� M� �� �t �� �t �� M�      3    , �� C� �h C� �h f� �� f� �� C�      3    , T� "�D `` "�D `` #�( T� #�( T� "�D      3    , `� !�� l< !�� l< "�� `� "�� `� !��      3    , o0 �P i0 �P i0 � o0 � o0 �P +  ,VR_NO_BUS       3    , .UT � .a � .a �� .UT �� .UT �      3    , 	�0 
�P 	�� 
�P 	�� � 	�0 � 	�0 
�P      3    , 4 �� %� �� %� 0  4 0  4 ��      3    , �� � �H � �H 0  �� 0  �� �      3    , %�� 	u� %�X 	u� %�X 	� %�� 	� %�� 	u�      3    , ![ %�L !f� %�L !f� %�t ![ %�t ![ %�L      3    ,  zt %�L  �, %�L  �, %�t  zt %�t  zt %�L      1    , 0
� � 0� � 0� � 0
� � 0
� �      1    , +]� \� ,� \� ,� hX +]� hX +]� \�      1    , -�| L� .2, L� .2, Xl -�| Xl -�| L�      1    , "�� H +�� H +�� #  "�� #  "�� H      1    , �� _D Kt _D Kt j� �� j� �� _D      1    , �� *h q@ *h q@ 6  �� 6  �� *h      1    , e$ z� �� z� �� �t e$ �t e$ z�      1    , ,� �� "� �� "� �8 ,� �8 ,� ��      1    , ut !, �T !, �T ,� ut ,� ut !,      1    , � H 
P� H 
P� #  � #  � H      1    , !�� \� "� \� "� hX !�� hX !�� \�      1    , !� � !�� � !�� �� !� �� !� �      1    , �� 
�P �� 
�P �� 
� �� 
� �� 
�P      1    , U� � $l8 � $l8 �� U� �� U� �      1    , !� �L "1� �L "1� � !� � !� �L      1    , wh �  �H �  �H �� wh �� wh �       1    , &�� 
�P *�� 
�P *�� 
� &�� 
� &�� 
�P      1    , !�P � ";� � ";� �� !�P �� !�P �      1    , Z� � �d � �d �� Z� �� Z� �      1    , q� �� ' �� ' �8 q� �8 q� ��      1    ,  �  C� �  C� ��  ��  �       1    , \x *h �L *h �L 6  \x 6  \x *h      1    , �H 6� \� 6� \� B@ �H B@ �H 6�      1    , )�� \� *!( \� *!( hX )�� hX )�� \�      1    , ,$� _D ,S� _D ,S� j� ,$� j� ,$� _D      1    , +d  Ĭ +@D  Ĭ +@D  �d +d  �d +d  Ĭ      1    , #�� 
�P $T� 
�P $T� 
� #�� 
� #�� 
�P      1    , �� �� �x �� �x �� �� �� �� ��      1    , -� �  .(h �  .(h �� -� �� -� �       1    ,  � f� �� f� �� r�  � r�  � f�      1    , *�p .P *�P .P *�P : *�p : *�p .P      1    , .� � ]� � ]� X .� X .� �      1    , �� � t � t %\ �� %\ �� �      1    , �$ �d O� �d O�  �$  �$ �d      1    , !� W� "5� W� "5� ct !� ct !� W�      1    , 	�  � 	�  � 	�  �� 	�  �� 	�  �      1    , � \� � \� � hX � hX � \�      1    ,  �D \�  �$ \�  �$ hX  �D hX  �D \�      1    , 	�4 U �L U �L `� 	�4 `� 	�4 U      1    , o� �� �` �� �` �� o� �� o� ��      1    , D M� q@ M� q@ YH D YH D M�      1    , �� H �L H �L #  �� #  �� H      1    , *@ ( *L  ( *L  � *@ � *@ (      1    , � _D �T _D �T j� � j� � _D      1    , �� _D iP _D iP j� �� j� �� _D      1    , !�  Ĭ !zP  Ĭ !zP  �d !�  �d !�  Ĭ      1    , �   Ĭ �   Ĭ �   �d �   �d �   Ĭ      1    , !�  �� !E�  �� !E�  � !�  � !�  ��      1    , Y� H _@ H _@ #  Y� #  Y� H      1    , �t Ӝ :� Ӝ :� �T �t �T �t Ӝ      1    , J �  x� �  x� �� J �� J �       1    , � �@ %y� �@ %y� �� � �� � �@      1    , "� Ӝ  p� Ӝ  p� �T "� �T "� Ӝ      1    , *�� ( +� ( +� � *�� � *�� (      1    , ,�h �  -�\ �  -�\ �� ,�h �� ,�h �       1    , ]0 �� ( �� ( �� ]0 �� ]0 ��      1    , ۴ Ӝ �  Ӝ �  �T ۴ �T ۴ Ӝ      1    , xd \� &8 \� &8 hX xd hX xd \�      1    , 24 � a � a �� 24 �� 24 �      1    , l  Ĭ �@  Ĭ �@  �d l  �d l  Ĭ      1    , g� $�� h $�� h %� g� %� g� $��      1    , �, [|  �� [|  �� g4 �, g4 �, [|      1    , �D !, h !, h ,� �D ,� �D !,      1    , o0 &�� Q� &�� Q� &�� o0 &�� o0 &�� +  ,VR_NO_BUS       1    , �� �$ �$ �$ �$ �� �� �� �� �$      1    , 
�� \� �� \� �� hX 
�� hX 
�� \�      1    , -p %$ 0rX %$ 0rX %=4 -p %=4 -p %$ +  ,VR_NO_BUS       1    , �< H &8 H &8 #  �< #  �< H      1    , ,x !, [X !, [X ,� ,x ,� ,x !,      1    , ( �  V� �  V� �� ( �� ( �       1    , $)� ~� $�� ~� $�� �< $)� �< $)� ~�      1    , Ĵ Ӝ � Ӝ � �T Ĵ �T Ĵ Ӝ      1    , )�  Ĭ )��  Ĭ )��  �d )�  �d )�  Ĭ      1    , _� _D �, _D �, j� _� j� _� _D      1    , @ ( �@ ( �@ � @ � @ (      1    , �� [| l` [| l` g4 �� g4 �� [|      1    , �$ *h �� *h �� 6  �$ 6  �$ *h      1    , �� �� � �� � �� �� �� �� ��      1    , v� � �� � �� �� v� �� v� �      1    , &�l 6� 'H 6� 'H B@ &�l B@ &�l 6�      1    , �t �d �D �d �D  �t  �t �d      1    , P � ]� � ]� �� P �� P �      1    , ( [| 4 [| 4 g4 ( g4 ( [|      1    , -p &�� /�h &�� /�h &�� -p &�� -p &�� +  ,VR_NO_BUS       1    , �� !, �H !, �H ,� �� ,� �� !,      1    , � ( � ( � � � � � (      1    , �� �  | �  | �� �� �� �� �       1    , �� Ӝ &� Ӝ &� �T �� �T �� Ӝ      1    , $P� 
�x $� 
�x $� 
�0 $P� 
�0 $P� 
�x      1    , `� Ӝ � Ӝ � �T `� �T `� Ӝ      1    ,  �@ %$ Q� %$ Q� %=4  �@ %=4  �@ %$ +  ,VR_NO_BUS       1    ,  �� %$  �@ %$  �@ %=4  �� %=4  �� %$ +  ,VR_NO_BUS       1    , !�X %$ !�@ %$ !�@ %=4 !�X %=4 !�X %$ +  ,VR_NO_BUS       1    , "1� %$ "M@ %$ "M@ %=4 "1� %=4 "1� %$ +  ,VR_NO_BUS       1    , #< %$ #(  %$ #(  %=4 #< %=4 #< %$ +  ,VR_NO_BUS       1    , %�� %$ &  %$ &  %=4 %�� %=4 %�� %$ +  ,VR_NO_BUS       1    , (� %$ )#@ %$ )#@ %=4 (� %=4 (� %$ +  ,VR_NO_BUS       1    , )� &�� )�  &�� )�  &�� )� &�� )� &�� +  ,VR_NO_BUS       1    , )� %$ )�  %$ )�  %=4 )� %=4 )� %$ +  ,VR_NO_BUS       1    , 	�0 
�P 
\X 
�P 
\X 
� 	�0 
� 	�0 
�P      1    , �� 
�P �d 
�P �d 
� �� 
� �� 
�P      1    , b� 
�P ! 
�P ! 
� b� 
� b� 
�P      1    , �� �  �@ �  �@ �� �� �� �� �       1    , #� 6� #�� 6� #�� B@ #� B@ #� 6�      1    , _� H �h H �h #  _� #  _� H      1    , �| _D %�( _D %�( j� �| j� �| _D      1    ,  | %$ *@ %$ *@ %=4  | %=4  | %$ +  ,VR_NO_BUS       1    ,  X %$ $@ %$ $@ %=4  X %=4  X %$ +  ,VR_NO_BUS       1    , X %$ @ %$ @ %=4 X %=4 X %$ +  ,VR_NO_BUS       1    , X %$ @ %$ @ %=4 X %=4 X %$ +  ,VR_NO_BUS       1    , �< %$ �  %$ �  %=4 �< %=4 �< %$ +  ,VR_NO_BUS       1    , � %$ �  %$ �  %=4 � %=4 � %$ +  ,VR_NO_BUS       1    , � %$ �  %$ �  %=4 � %=4 � %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , [| %$ e@ %$ e@ %=4 [| %=4 [| %$ +  ,VR_NO_BUS       1    , [X %$ _@ %$ _@ %=4 [X %=4 [X %$ +  ,VR_NO_BUS       1    ,  UX %$  Y@ %$  Y@ %=4  UX %=4  UX %$ +  ,VR_NO_BUS       1    , �h %$ �� %$ �� %=4 �h %=4 �h %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , 	h %$ 	'� %$ 	'� %=4 	h %=4 	h %$ +  ,VR_NO_BUS       1    , 
� %$ 
!� %$ 
!� %=4 
� %=4 
� %$ +  ,VR_NO_BUS       1    , 
�� %$ 
�  %$ 
�  %=4 
�� %=4 
�� %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , ,� %$ H@ %$ H@ %=4 ,� %=4 ,� %$ +  ,VR_NO_BUS       1    , �h %$ � %$ � %=4 �h %=4 �h %$ +  ,VR_NO_BUS       1    , Լ %$ ހ %$ ހ %=4 Լ %=4 Լ %$ +  ,VR_NO_BUS       1    , Ԙ %$ ؀ %$ ؀ %=4 Ԙ %=4 Ԙ %$ +  ,VR_NO_BUS       1    , :( %$ U� %$ U� %=4 :( %=4 :( %$ +  ,VR_NO_BUS       1    , K� %$ O� %$ O� %=4 K� %=4 K� %$ +  ,VR_NO_BUS       1    , #� #� #�  #� #�  #5� #� #5� #� #� +  ,VR_NO_BUS       1    , $u� #� $� #� $� #5� $u� #5� $u� #� +  ,VR_NO_BUS       1    , %u� #� %y� #� %y� #5� %u� #5� %u� #� +  ,VR_NO_BUS       1    , &J� #� &T� #� &T� #5� &J� #5� &J� #� +  ,VR_NO_BUS       1    , 'J� #� 'N� #� 'N� #5� 'J� #5� 'J� #� +  ,VR_NO_BUS       1    , *!( #� *<� #� *<� #5� *!( #5� *!( #� +  ,VR_NO_BUS       1    , -( #� -*� #� -*� #5� -( #5� -( #� +  ,VR_NO_BUS       1    , -̜ #� -�  #� -�  #5� -̜ #5� -̜ #� +  ,VR_NO_BUS       1    , .�( #� 0rX #� 0rX #5� .�( #5� .�( #� +  ,VR_NO_BUS       1    ,  �@ #� Q� #� Q� #5�  �@ #5�  �@ #� +  ,VR_NO_BUS       1    , �� %$ @ %$ @ %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , �h %$ �� %$ �� %=4 �h %=4 �h %$ +  ,VR_NO_BUS       1    , �� %$ �� %$ �� %=4 �� %=4 �� %$ +  ,VR_NO_BUS       1    , C� %$ _  %$ _  %=4 C� %=4 C� %$ +  ,VR_NO_BUS       1    , /� %$ 9� %$ 9� %=4 /� %=4 /� %$ +  ,VR_NO_BUS       1    , X #� @ #� @ #5� X #5� X #� +  ,VR_NO_BUS       1    , y� #� �@ #� �@ #5� y� #5� y� #� +  ,VR_NO_BUS       1    , s� #� �@ #� �@ #5� s� #5� s� #� +  ,VR_NO_BUS       1    , `< #� j  #� j  #5� `< #5� `< #� +  ,VR_NO_BUS       1    , ` #� d  #� d  #5� ` #5� ` #� +  ,VR_NO_BUS       1    , 4� #� >� #� >� #5� 4� #5� 4� #� +  ,VR_NO_BUS       1    , 4� #� 8� #� 8� #5� 4� #5� 4� #� +  ,VR_NO_BUS       1    , .� #� 2� #� 2� #5� .� #5� .� #� +  ,VR_NO_BUS       1    , (� #� ,� #� ,� #5� (� #5� (� #� +  ,VR_NO_BUS       1    , �� #� � #� � #5� �� #5� �� #� +  ,VR_NO_BUS       1    , �� #� � #� � #5� �� #5� �� #� +  ,VR_NO_BUS       1    , �| #� �@ #� �@ #5� �| #5� �| #� +  ,VR_NO_BUS       1    ,  �< #�  �  #�  �  #5�  �< #5�  �< #� +  ,VR_NO_BUS       1    , !� #� !�  #� !�  #5� !� #5� !� #� +  ,VR_NO_BUS       1    , "� #� "�  #� "�  #5� "� #5� "� #� +  ,VR_NO_BUS       1    , �| #� �@ #� �@ #5� �| #5� �| #� +  ,VR_NO_BUS       1    , 	�X #� 	�@ #� 	�@ #5� 	�X #5� 	�X #� +  ,VR_NO_BUS       1    , 
�X #� 
�@ #� 
�@ #5� 
�X #5� 
�X #� +  ,VR_NO_BUS       1    , �X #� �@ #� �@ #5� �X #5� �X #� +  ,VR_NO_BUS       1    , �X #� �@ #� �@ #5� �X #5� �X #� +  ,VR_NO_BUS       1    , �< #� �  #� �  #5� �< #5� �< #� +  ,VR_NO_BUS       1    , � #� �  #� �  #5� � #5� � #� +  ,VR_NO_BUS       1    , � #� #  #� #  #5� � #5� � #� +  ,VR_NO_BUS       1    ,  #�   #�   #5�  #5�  #� +  ,VR_NO_BUS       1    , �� #� �� #� �� #5� �� #5� �� #� +  ,VR_NO_BUS       1    , �� #� �� #� �� #5� �� #5� �� #� +  ,VR_NO_BUS       1    , Sh #� n� #� n� #5� Sh #5� Sh #� +  ,VR_NO_BUS       1    , d� #� h� #� h� #5� d� #5� d� #� +  ,VR_NO_BUS       1    , 9� #� C� #� C� #5� 9� #5� 9� #� +  ,VR_NO_BUS       1    , | #� @ #� @ #5� | #5� | #� +  ,VR_NO_BUS       1    , (�X ! (�@ ! (�@ !.$ (�X !.$ (�X ! +  ,VR_NO_BUS       1    , )w< ! )�  ! )�  !.$ )w< !.$ )w< ! +  ,VR_NO_BUS       1    , )� ! )�  ! )�  !.$ )� !.$ )� ! +  ,VR_NO_BUS       1    , *� ! *�  ! *�  !.$ *� !.$ *� ! +  ,VR_NO_BUS       1    , +�� ! +�� ! +�� !.$ +�� !.$ +�� ! +  ,VR_NO_BUS       1    , ,�� ! ,�� ! ,�� !.$ ,�� !.$ ,�� ! +  ,VR_NO_BUS       1    , -�� ! 0rX ! 0rX !.$ -�� !.$ -�� ! +  ,VR_NO_BUS       1    ,  �@ ! Q� ! Q� !.$  �@ !.$  �@ ! +  ,VR_NO_BUS       1    , Ҩ #� �  #� �  #5� Ҩ #5� Ҩ #� +  ,VR_NO_BUS       1    , � #� �  #� �  #5� � #5� � #� +  ,VR_NO_BUS       1    , I� #� e  #� e  #5� I� #5� I� #� +  ,VR_NO_BUS       1    , 5� #� ?� #� ?� #5� 5� #5� 5� #� +  ,VR_NO_BUS       1    , 5� #� 9� #� 9� #5� 5� #5� 5� #� +  ,VR_NO_BUS       1    , /� #� 3� #� 3� #5� /� #5� /� #� +  ,VR_NO_BUS       1    , � #� � #� � #5� � #5� � #� +  ,VR_NO_BUS       1    , h ! 8� ! 8� !.$ h !.$ h ! +  ,VR_NO_BUS       1    , .� ! 2� ! 2� !.$ .� !.$ .� ! +  ,VR_NO_BUS       1    , � ! � ! � !.$ � !.$ � ! +  ,VR_NO_BUS       1    , � ! � ! � !.$ � !.$ � ! +  ,VR_NO_BUS       1    , �� ! � ! � !.$ �� !.$ �� ! +  ,VR_NO_BUS       1    , �| ! �@ ! �@ !.$ �| !.$ �| ! +  ,VR_NO_BUS       1    ,  �X !  �@ !  �@ !.$  �X !.$  �X ! +  ,VR_NO_BUS       1    , !�< ! !�  ! !�  !.$ !�< !.$ !�< ! +  ,VR_NO_BUS       1    , "� ! "�  ! "�  !.$ "� !.$ "� ! +  ,VR_NO_BUS       1    , #{� ! #�� ! #�� !.$ #{� !.$ #{� ! +  ,VR_NO_BUS       1    , $V� ! $`� ! $`� !.$ $V� !.$ $V� ! +  ,VR_NO_BUS       1    , %V� ! %Z� ! %Z� !.$ %V� !.$ %V� ! +  ,VR_NO_BUS       1    , &+| ! &5@ ! &5@ !.$ &+| !.$ &+| ! +  ,VR_NO_BUS       1    , &�� ! &�@ ! &�@ !.$ &�� !.$ &�� ! +  ,VR_NO_BUS       1    , '�X ! '�@ ! '�@ !.$ '�X !.$ '�X ! +  ,VR_NO_BUS       1    , ژ ! ހ ! ހ !.$ ژ !.$ ژ ! +  ,VR_NO_BUS       1    , _h ! z� ! z� !.$ _h !.$ _h ! +  ,VR_NO_BUS       1    , � ! 6@ ! 6@ !.$ � !.$ � ! +  ,VR_NO_BUS       1    , �h ! �� ! �� !.$ �h !.$ �h ! +  ,VR_NO_BUS       1    , Sh ! n� ! n� !.$ Sh !.$ Sh ! +  ,VR_NO_BUS       1    , ?� ! I� ! I� !.$ ?� !.$ ?� ! +  ,VR_NO_BUS       1    , | ! $@ ! $@ !.$ | !.$ | ! +  ,VR_NO_BUS       1    , X ! @ ! @ !.$ X !.$ X ! +  ,VR_NO_BUS       1    , X ! @ ! @ !.$ X !.$ X ! +  ,VR_NO_BUS       1    , y� ! �@ ! �@ !.$ y� !.$ y� ! +  ,VR_NO_BUS       1    , f< ! p  ! p  !.$ f< !.$ f< ! +  ,VR_NO_BUS       1    , Ѩ ! �  ! �  !.$ Ѩ !.$ Ѩ ! +  ,VR_NO_BUS       1    , � ! �  ! �  !.$ � !.$ � ! +  ,VR_NO_BUS       1    , � ! �  ! �  !.$ � !.$ � ! +  ,VR_NO_BUS       1    , �� ! �� ! �� !.$ �� !.$ �� ! +  ,VR_NO_BUS       1    , G� ! K� ! K� !.$ G� !.$ G� ! +  ,VR_NO_BUS       1    , �� ! @ ! @ !.$ �� !.$ �� ! +  ,VR_NO_BUS       1    , �h ! �� ! �� !.$ �h !.$ �h ! +  ,VR_NO_BUS       1    , �� ! �� ! �� !.$ �� !.$ �� ! +  ,VR_NO_BUS       1    , �� ! �� ! �� !.$ �� !.$ �� ! +  ,VR_NO_BUS       1    , h ! 3� ! 3� !.$ h !.$ h ! +  ,VR_NO_BUS       1    , )� ! -� ! -� !.$ )� !.$ )� ! +  ,VR_NO_BUS       1    , 	#� ! 	'� ! 	'� !.$ 	#� !.$ 	#� ! +  ,VR_NO_BUS       1    , 	�� ! 
� ! 
� !.$ 	�� !.$ 	�� ! +  ,VR_NO_BUS       1    , 
�� ! 
�� ! 
�� !.$ 
�� !.$ 
�� ! +  ,VR_NO_BUS       1    , � ! �� ! �� !.$ � !.$ � ! +  ,VR_NO_BUS       1    , wh ! �� ! �� !.$ wh !.$ wh ! +  ,VR_NO_BUS       1    , c� ! m� ! m� !.$ c� !.$ c� ! +  ,VR_NO_BUS       1    , �( ! � ! � !.$ �( !.$ �( ! +  ,VR_NO_BUS       1    , �� ! � ! � !.$ �� !.$ �� ! +  ,VR_NO_BUS       1    , #$ �d #(  �d #(  t #$ t #$ �d +  ,VR_NO_BUS       1    , #�� �d $� �d $� t #�� t #�� �d +  ,VR_NO_BUS       1    , $�� �d $�� �d $�� t $�� t $�� �d +  ,VR_NO_BUS       1    , %�� �d %�� �d %�� t %�� t %�� �d +  ,VR_NO_BUS       1    , &Ǽ �d &р �d &р t &Ǽ t &Ǽ �d +  ,VR_NO_BUS       1    , 'ǘ �d 'ˀ �d 'ˀ t 'ǘ t 'ǘ �d +  ,VR_NO_BUS       1    , (�| �d (�@ �d (�@ t (�| t (�| �d +  ,VR_NO_BUS       1    , )�X �d )�@ �d )�@ t )�X t )�X �d +  ,VR_NO_BUS       1    , *q< �d *{  �d *{  t *q< t *q< �d +  ,VR_NO_BUS       1    , +q �d +u  �d +u  t +q t +q �d +  ,VR_NO_BUS       1    , ,k �d ,o  �d ,o  t ,k t ,k �d +  ,VR_NO_BUS       1    , -?� �d -I� �d -I� t -?� t -?� �d +  ,VR_NO_BUS       1    , .� �d .$� �d .$� t .� t .� �d +  ,VR_NO_BUS       1    , .�( �d 0rX �d 0rX t .�( t .�( �d +  ,VR_NO_BUS       1    ,  �@ �d Q� �d Q� t  �@ t  �@ �d +  ,VR_NO_BUS       1    , r< �d |  �d |  t r< t r< �d +  ,VR_NO_BUS       1    , r �d v  �d v  t r t r �d +  ,VR_NO_BUS       1    , l �d p  �d p  t l t l �d +  ,VR_NO_BUS       1    , @� �d J� �d J� t @� t @� �d +  ,VR_NO_BUS       1    , @� �d D� �d D� t @� t @� �d +  ,VR_NO_BUS       1    , :� �d >� �d >� t :� t :� �d +  ,VR_NO_BUS       1    , � �d � �d � t � t � �d +  ,VR_NO_BUS       1    , � �d � �d � t � t � �d +  ,VR_NO_BUS       1    , 	� �d � �d � t 	� t 	� �d +  ,VR_NO_BUS       1    , o( �d �� �d �� t o( t o( �d +  ,VR_NO_BUS       1    , [| �d e@ �d e@ t [| t [| �d +  ,VR_NO_BUS       1    , [X �d _@ �d _@ t [X t [X �d +  ,VR_NO_BUS       1    ,  0< �d  :  �d  :  t  0< t  0< �d +  ,VR_NO_BUS       1    , !0 �d !4  �d !4  t !0 t !0 �d +  ,VR_NO_BUS       1    , "* �d ".  �d ".  t "* t "* �d +  ,VR_NO_BUS       1    , �� �d �� �d �� t �� t �� �d +  ,VR_NO_BUS       1    , 	�� �d 	�� �d 	�� t 	�� t 	�� �d +  ,VR_NO_BUS       1    , 
{� �d 
� �d 
� t 
{� t 
{� �d +  ,VR_NO_BUS       1    , u� �d y� �d y� t u� t u� �d +  ,VR_NO_BUS       1    , � �d 5  �d 5  t � t � �d +  ,VR_NO_BUS       1    , + �d /  �d /  t + t + �d +  ,VR_NO_BUS       1    , �( �d � �d � t �( t �( �d +  ,VR_NO_BUS       1    , �� �d � �d � t �� t �� �d +  ,VR_NO_BUS       1    , �| �d �@ �d �@ t �| t �| �d +  ,VR_NO_BUS       1    , �X �d �@ �d �@ t �X t �X �d +  ,VR_NO_BUS       1    , �< �d �  �d �  t �< t �< �d +  ,VR_NO_BUS       1    , � �d �  �d �  t � t � �d +  ,VR_NO_BUS       1    , � �d *@ �d *@ t � t � �d +  ,VR_NO_BUS       1    , �� �d �@ �d �@ t �� t �� �d +  ,VR_NO_BUS       1    , �X �d �@ �d �@ t �X t �X �d +  ,VR_NO_BUS       1    , (%X s4 ()@ s4 ()@ �D (%X �D (%X s4 +  ,VR_NO_BUS       1    , )X s4 )#@ s4 )#@ �D )X �D )X s4 +  ,VR_NO_BUS       1    , )�< s4 )�  s4 )�  �D )�< �D )�< s4 +  ,VR_NO_BUS       1    , *� s4 *�  s4 *�  �D *� �D *� s4 +  ,VR_NO_BUS       1    , +�� s4 +�� s4 +�� �D +�� �D +�� s4 +  ,VR_NO_BUS       1    , ,�� s4 ,�� s4 ,�� �D ,�� �D ,�� s4 +  ,VR_NO_BUS       1    , -�� s4 -�� s4 -�� �D -�� �D -�� s4 +  ,VR_NO_BUS       1    , .�� s4 0rX s4 0rX �D .�� �D .�� s4 +  ,VR_NO_BUS       1    ,  �@ s4 Q� s4 Q� �D  �@ �D  �@ s4 +  ,VR_NO_BUS       1    , G� �d K� �d K� t G� t G� �d +  ,VR_NO_BUS       1    , �h �d �� �d �� t �h t �h �d +  ,VR_NO_BUS       1    , �� �d �� �d �� t �� t �� �d +  ,VR_NO_BUS       1    , �� �d �� �d �� t �� t �� �d +  ,VR_NO_BUS       1    , �� �d �� �d �� t �� t �� �d +  ,VR_NO_BUS       1    , �� �d �� �d �� t �� t �� �d +  ,VR_NO_BUS       1    , �( s4 �� s4 �� �D �( �D �( s4 +  ,VR_NO_BUS       1    , �� s4 �� s4 �� �D �� �D �� s4 +  ,VR_NO_BUS       1    , �� s4 �� s4 �� �D �� �D �� s4 +  ,VR_NO_BUS       1    , a| s4 k@ s4 k@ �D a| �D a| s4 +  ,VR_NO_BUS       1    , aX s4 e@ s4 e@ �D aX �D aX s4 +  ,VR_NO_BUS       1    , [X s4 _@ s4 _@ �D [X �D [X s4 +  ,VR_NO_BUS       1    , �� s4 �@ s4 �@ �D �� �D �� s4 +  ,VR_NO_BUS       1    ,  �X s4  �@ s4  �@ �D  �X �D  �X s4 +  ,VR_NO_BUS       1    , !�< s4 !�  s4 !�  �D !�< �D !�< s4 +  ,VR_NO_BUS       1    , "�� s4 "�� s4 "�� �D "�� �D "�� s4 +  ,VR_NO_BUS       1    , #�� s4 #�� s4 #�� �D #�� �D #�� s4 +  ,VR_NO_BUS       1    , ${� s4 $� s4 $� �D ${� �D ${� s4 +  ,VR_NO_BUS       1    , %P� s4 %Z� s4 %Z� �D %P� �D %P� s4 +  ,VR_NO_BUS       1    , &P� s4 &T� s4 &T� �D &P� �D &P� s4 +  ,VR_NO_BUS       1    , '%| s4 '/@ s4 '/@ �D '%| �D '%| s4 +  ,VR_NO_BUS       1    , � s4 � s4 � �D � �D � s4 +  ,VR_NO_BUS       1    , �� s4 � s4 � �D �� �D �� s4 +  ,VR_NO_BUS       1    , �| s4 �@ s4 �@ �D �| �D �| s4 +  ,VR_NO_BUS       1    , �X s4 �@ s4 �@ �D �X �D �X s4 +  ,VR_NO_BUS       1    , � s4 6@ s4 6@ �D � �D � s4 +  ,VR_NO_BUS       1    , ,X s4 0@ s4 0@ �D ,X �D ,X s4 +  ,VR_NO_BUS       1    , &X s4 *@ s4 *@ �D &X �D &X s4 +  ,VR_NO_BUS       1    ,  X s4 $@ s4 $@ �D  X �D  X s4 +  ,VR_NO_BUS       1    , �< s4 �  s4 �  �D �< �D �< s4 +  ,VR_NO_BUS       1    , � s4 �  s4 �  �D � �D � s4 +  ,VR_NO_BUS       1    , �� s4 �� s4 �� �D �� �D �� s4 +  ,VR_NO_BUS       1    , 5h s4 P� s4 P� �D 5h �D 5h s4 +  ,VR_NO_BUS       1    , F� s4 J� s4 J� �D F� �D F� s4 +  ,VR_NO_BUS       1    , @� s4 D� s4 D� �D @� �D @� s4 +  ,VR_NO_BUS       1    , � s4 � s4 � �D � �D � s4 +  ,VR_NO_BUS       1    , .�� 8� 0rX 8� 0rX _� .�� _� .�� 8� +  ,VR_NO_BUS       1    ,  �@ 8� Q� 8� Q� _�  �@ _�  �@ 8� +  ,VR_NO_BUS       1    , �h s4 �� s4 �� �D �h �D �h s4 +  ,VR_NO_BUS       1    , �� s4 �� s4 �� �D �� �D �� s4 +  ,VR_NO_BUS       1    , �� s4 �� s4 �� �D �� �D �� s4 +  ,VR_NO_BUS       1    , C� s4 _  s4 _  �D C� �D C� s4 +  ,VR_NO_BUS       1    , U s4 Y  s4 Y  �D U �D U s4 +  ,VR_NO_BUS       1    , �( s4 � s4 � �D �( �D �( s4 +  ,VR_NO_BUS       1    , �� s4 �  s4 �  �D �� �D �� s4 +  ,VR_NO_BUS       1    , � s4 �  s4 �  �D � �D � s4 +  ,VR_NO_BUS       1    , 	�� s4 	�� s4 	�� �D 	�� �D 	�� s4 +  ,VR_NO_BUS       1    , 
�� s4 
�� s4 
�� �D 
�� �D 
�� s4 +  ,VR_NO_BUS       1    , o� s4 y� s4 y� �D o� �D o� s4 +  ,VR_NO_BUS       1    , o� s4 s� s4 s� �D o� �D o� s4 +  ,VR_NO_BUS       1    , �( s4 �� s4 �� �D �( �D �( s4 +  ,VR_NO_BUS       1    , !� 8� !� 8� !� _� !� _� !� 8� +  ,VR_NO_BUS       1    , "� 8� "� 8� "� _� "� _� "� 8� +  ,VR_NO_BUS       1    , #ߘ 8� #� 8� #� _� #ߘ _� #ߘ 8� +  ,VR_NO_BUS       1    , $E( 8� $`� 8� $`� _� $E( _� $E( 8� +  ,VR_NO_BUS       1    , %1| 8� %;@ 8� %;@ _� %1| _� %1| 8� +  ,VR_NO_BUS       1    , &1X 8� &5@ 8� &5@ _� &1X _� &1X 8� +  ,VR_NO_BUS       1    , '+X 8� '/@ 8� '/@ _� '+X _� '+X 8� +  ,VR_NO_BUS       1    , '� 8� (
  8� (
  _� '� _� '� 8� +  ,VR_NO_BUS       1    , (k� 8� (�  8� (�  _� (k� _� (k� 8� +  ,VR_NO_BUS       1    , )} 8� )�  8� )�  _� )} _� )} 8� +  ,VR_NO_BUS       1    , *w 8� *{  8� *{  _� *w _� *w 8� +  ,VR_NO_BUS       1    , +K� 8� +U� 8� +U� _� +K� _� +K� 8� +  ,VR_NO_BUS       1    , ,K� 8� ,O� 8� ,O� _� ,K� _� ,K� 8� +  ,VR_NO_BUS       1    , - � 8� -*� 8� -*� _� - � _� - � 8� +  ,VR_NO_BUS       1    , -�( 8� -�� 8� -�� _� -�( _� -�( 8� +  ,VR_NO_BUS       1    , f� 8� �  8� �  _� f� _� f� 8� +  ,VR_NO_BUS       1    , R� 8� \� 8� \� _� R� _� R� 8� +  ,VR_NO_BUS       1    , R� 8� V� 8� V� _� R� _� R� 8� +  ,VR_NO_BUS       1    , L� 8� P� 8� P� _� L� _� L� 8� +  ,VR_NO_BUS       1    , !� 8� +� 8� +� _� !� _� !� 8� +  ,VR_NO_BUS       1    , !� 8� %� 8� %� _� !� _� !� 8� +  ,VR_NO_BUS       1    , � 8� � 8� � _� � _� � 8� +  ,VR_NO_BUS       1    , �| 8� �@ 8� �@ _� �| _� �| 8� +  ,VR_NO_BUS       1    , [� 8� w@ 8� w@ _� [� _� [� 8� +  ,VR_NO_BUS       1    , H< 8� R  8� R  _� H< _� H< 8� +  ,VR_NO_BUS       1    , H 8� L  8� L  _� H _� H 8� +  ,VR_NO_BUS       1    , B 8� F  8� F  _� B _� B 8� +  ,VR_NO_BUS       1    , � 8�  � 8�  � _� � _� � 8� +  ,VR_NO_BUS       1    , � 8� �� 8� �� _� � _� � 8� +  ,VR_NO_BUS       1    ,  � 8�  �� 8�  �� _�  � _�  � 8� +  ,VR_NO_BUS       1    , �� 8� �� 8� �� _� �� _� �� 8� +  ,VR_NO_BUS       1    , 	h 8� 	'� 8� 	'� _� 	h _� 	h 8� +  ,VR_NO_BUS       1    , 	�� 8� 
� 8� 
� _� 	�� _� 	�� 8� +  ,VR_NO_BUS       1    , 
�� 8� 
�� 8� 
�� _� 
�� _� 
�� 8� +  ,VR_NO_BUS       1    , ^( 8� y� 8� y� _� ^( _� ^( 8� +  ,VR_NO_BUS       1    , J| 8� T@ 8� T@ _� J| _� J| 8� +  ,VR_NO_BUS       1    , %< 8� /  8� /  _� %< _� %< 8� +  ,VR_NO_BUS       1    , % 8� )  8� )  _� % _� % 8� +  ,VR_NO_BUS       1    , �� 8� � 8� � _� �� _� �� 8� +  ,VR_NO_BUS       1    , �� 8� �� 8� �� _� �� _� �� 8� +  ,VR_NO_BUS       1    , �� 8� �@ 8� �@ _� �� _� �� 8� +  ,VR_NO_BUS       1    , �X 8� �@ 8� �@ _� �X _� �X 8� +  ,VR_NO_BUS       1    , �< 8� �  8� �  _� �< _� �< 8� +  ,VR_NO_BUS       1    , � 8�   8�   _� � _� � 8� +  ,VR_NO_BUS       1    ,  8�   8�   _�  _�  8� +  ,VR_NO_BUS       1    , 'ǘ  'ˀ  'ˀ 9, 'ǘ 9, 'ǘ  +  ,VR_NO_BUS       1    , (��  (ŀ  (ŀ 9, (�� 9, (��  +  ,VR_NO_BUS       1    , )�|  )�@  )�@ 9, )�| 9, )�|  +  ,VR_NO_BUS       1    , *�X  *�@  *�@ 9, *�X 9, *�X  +  ,VR_NO_BUS       1    , +�X  +�@  +�@ 9, +�X 9, +�X  +  ,VR_NO_BUS       1    , ,S�  ,o   ,o  9, ,S� 9, ,S�  +  ,VR_NO_BUS       1    , -e  -i   -i  9, -e 9, -e  +  ,VR_NO_BUS       1    , -ʨ  0rX  0rX 9, -ʨ 9, -ʨ  +  ,VR_NO_BUS       1    ,  �@  Q�  Q� 9,  �@ 9,  �@  +  ,VR_NO_BUS       1    , "� 8� ,� 8� ,� _� "� _� "� 8� +  ,VR_NO_BUS       1    , "� 8� &� 8� &� _� "� _� "� 8� +  ,VR_NO_BUS       1    , � 8�  � 8�  � _� � _� � 8� +  ,VR_NO_BUS       1    , �� 8� �  8� �  _� �� _� �� 8� +  ,VR_NO_BUS       1    , �� 8� �� 8� �� _� �� _� �� 8� +  ,VR_NO_BUS       1    , �� 8� �� 8� �� _� �� _� �� 8� +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , g|  q@  q@ 9, g| 9, g|  +  ,VR_NO_BUS       1    , gX  k@  k@ 9, gX 9, gX  +  ,VR_NO_BUS       1    , aX  e@  e@ 9, aX 9, aX  +  ,VR_NO_BUS       1    , [X  _@  _@ 9, [X 9, [X  +  ,VR_NO_BUS       1    , ��  �@  �@ 9, �� 9, ��  +  ,VR_NO_BUS       1    ,  �X   �@   �@ 9,  �X 9,  �X  +  ,VR_NO_BUS       1    , !�<  !�   !�  9, !�< 9, !�<  +  ,VR_NO_BUS       1    , "�  "�   "�  9, "� 9, "�  +  ,VR_NO_BUS       1    , #{�  #��  #�� 9, #{� 9, #{�  +  ,VR_NO_BUS       1    , ${�  $�  $� 9, ${� 9, ${�  +  ,VR_NO_BUS       1    , %u�  %y�  %y� 9, %u� 9, %u�  +  ,VR_NO_BUS       1    , %�h  %��  %�� 9, %�h 9, %�h  +  ,VR_NO_BUS       1    , &Ǽ  &р  &р 9, &Ǽ 9, &Ǽ  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ]�  g�  g� 9, ]� 9, ]�  +  ,VR_NO_BUS       1    , ]�  a�  a� 9, ]� 9, ]�  +  ,VR_NO_BUS       1    , 2|  <@  <@ 9, 2| 9, 2|  +  ,VR_NO_BUS       1    , 2X  6@  6@ 9, 2X 9, 2X  +  ,VR_NO_BUS       1    , ,X  0@  0@ 9, ,X 9, ,X  +  ,VR_NO_BUS       1    , <       9, < 9, <  +  ,VR_NO_BUS       1    ,        9,  9,   +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , ,�h �T ,�� �T ,�� d ,�h d ,�h �T +  ,VR_NO_BUS       1    , -�h �T -�� �T -�� d -�h d -�h �T +  ,VR_NO_BUS       1    , .�� �T 0rX �T 0rX d .�� d .�� �T +  ,VR_NO_BUS       1    ,  �@ �T Q� �T Q� d  �@ d  �@ �T +  ,VR_NO_BUS       1    , G�  K�  K� 9, G� 9, G�  +  ,VR_NO_BUS       1    , ��  @  @ 9, �� 9, ��  +  ,VR_NO_BUS       1    , �X  @  @ 9, �X 9, �X  +  ,VR_NO_BUS       1    , �X  �@  �@ 9, �X 9, �X  +  ,VR_NO_BUS       1    , �<  �   �  9, �< 9, �<  +  ,VR_NO_BUS       1    , 7�  S   S  9, 7� 9, 7�  +  ,VR_NO_BUS       1    , I  M   M  9, I 9, I  +  ,VR_NO_BUS       1    , ��  �   �  9, �� 9, ��  +  ,VR_NO_BUS       1    , 	��  	��  	�� 9, 	�� 9, 	��  +  ,VR_NO_BUS       1    , 
��  
��  
�� 9, 
�� 9, 
��  +  ,VR_NO_BUS       1    , ��  ��  �� 9, �� 9, ��  +  ,VR_NO_BUS       1    , �X �T �@ �T �@ d �X d �X �T +  ,VR_NO_BUS       1    , �< �T �  �T �  d �< d �< �T +  ,VR_NO_BUS       1    ,  � �T  �  �T  �  d  � d  � �T +  ,VR_NO_BUS       1    , !� �T !�  �T !�  d !� d !� �T +  ,VR_NO_BUS       1    , "�� �T "�� �T "�� d "�� d "�� �T +  ,VR_NO_BUS       1    , #�� �T #�� �T #�� d #�� d #�� �T +  ,VR_NO_BUS       1    , ${� �T $� �T $� d ${� d ${� �T +  ,VR_NO_BUS       1    , %P� �T %Z� �T %Z� d %P� d %P� �T +  ,VR_NO_BUS       1    , &P� �T &T� �T &T� d &P� d &P� �T +  ,VR_NO_BUS       1    , 'J� �T 'N� �T 'N� d 'J� d 'J� �T +  ,VR_NO_BUS       1    , (| �T ()@ �T ()@ d (| d (| �T +  ,VR_NO_BUS       1    , )X �T )#@ �T )#@ d )X d )X �T +  ,VR_NO_BUS       1    , *X �T *@ �T *@ d *X d *X �T +  ,VR_NO_BUS       1    , *�< �T *�  �T *�  d *�< d *�< �T +  ,VR_NO_BUS       1    , +� �T ,O� �T ,O� d +� d +� �T +  ,VR_NO_BUS       1    , �h �T �� �T �� d �h d �h �T +  ,VR_NO_BUS       1    , ¼ �T ̀ �T ̀ d ¼ d ¼ �T +  ,VR_NO_BUS       1    ,  �T ƀ �T ƀ d  d  �T +  ,VR_NO_BUS       1    , (( �T C� �T C� d (( d (( �T +  ,VR_NO_BUS       1    , | �T @ �T @ d | d | �T +  ,VR_NO_BUS       1    , X �T @ �T @ d X d X �T +  ,VR_NO_BUS       1    , X �T @ �T @ d X d X �T +  ,VR_NO_BUS       1    , X �T @ �T @ d X d X �T +  ,VR_NO_BUS       1    , �< �T �  �T �  d �< d �< �T +  ,VR_NO_BUS       1    , �� �T �� �T �� d �� d �� �T +  ,VR_NO_BUS       1    , �� �T �� �T �� d �� d �� �T +  ,VR_NO_BUS       1    , �� �T �� �T �� d �� d �� �T +  ,VR_NO_BUS       1    , �( �T � �T � d �( d �( �T +  ,VR_NO_BUS       1    , �| �T �@ �T �@ d �| d �| �T +  ,VR_NO_BUS       1    , �X �T �@ �T �@ d �X d �X �T +  ,VR_NO_BUS       1    , � �T �  �T �  d � d � �T +  ,VR_NO_BUS       1    , �� �T �� �T �� d �� d �� �T +  ,VR_NO_BUS       1    , h �T -� �T -� d h d h �T +  ,VR_NO_BUS       1    , 	#� �T 	'� �T 	'� d 	#� d 	#� �T +  ,VR_NO_BUS       1    , 	�� �T 	�  �T 	�  d 	�� d 	�� �T +  ,VR_NO_BUS       1    , 
d( �T 
� �T 
� d 
d( d 
d( �T +  ,VR_NO_BUS       1    , P| �T Z@ �T Z@ d P| d P| �T +  ,VR_NO_BUS       1    , �� �T �@ �T �@ d �� d �� �T +  ,VR_NO_BUS       1    , 8� �T T@ �T T@ d 8� d 8� �T +  ,VR_NO_BUS       1    , %< �T /  �T /  d %< d %< �T +  ,VR_NO_BUS       1    , �� �T �  �T �  d �� d �� �T +  ,VR_NO_BUS       1    , � �T �  �T �  d � d � �T +  ,VR_NO_BUS       1    , � �T �  �T �  d � d � �T +  ,VR_NO_BUS       1    , � �T �  �T �  d � d � �T +  ,VR_NO_BUS       1    , j� �T t� �T t� d j� d j� �T +  ,VR_NO_BUS       1    , ( < Č (
  Č (
  � ( < � ( < Č +  ,VR_NO_BUS       1    , (�( Č (ŀ Č (ŀ � (�( � (�( Č +  ,VR_NO_BUS       1    , )�� Č )�� Č )�� � )�� � )�� Č +  ,VR_NO_BUS       1    , *@h Č *[� Č *[� � *@h � *@h Č +  ,VR_NO_BUS       1    , +Q� Č +U� Č +U� � +Q� � +Q� Č +  ,VR_NO_BUS       1    , ,&� Č ,0� Č ,0� � ,&� � ,&� Č +  ,VR_NO_BUS       1    , -&� Č -*� Č -*� � -&� � -&� Č +  ,VR_NO_BUS       1    , -ʨ Č -�  Č -�  � -ʨ � -ʨ Č +  ,VR_NO_BUS       1    , .f� Č 0rX Č 0rX � .f� � .f� Č +  ,VR_NO_BUS       1    ,  �@ Č Q� Č Q� �  �@ �  �@ Č +  ,VR_NO_BUS       1    , Ҩ �T �  �T �  d Ҩ d Ҩ �T +  ,VR_NO_BUS       1    , �( �T �� �T �� d �( d �( �T +  ,VR_NO_BUS       1    , �� �T �� �T �� d �� d �� �T +  ,VR_NO_BUS       1    , ( �T  � �T  � d ( d ( �T +  ,VR_NO_BUS       1    , �� �T �  �T �  d �� d �� �T +  ,VR_NO_BUS       1    , � Č �  Č �  � � � � Č +  ,VR_NO_BUS       1    , �� Č �� Č �� � �� � �� Č +  ,VR_NO_BUS       1    , �� Č �� Č �� � �� � �� Č +  ,VR_NO_BUS       1    , �� Č �� Č �� � �� � �� Č +  ,VR_NO_BUS       1    , z� Č �� Č �� � z� � z� Č +  ,VR_NO_BUS       1    , z� Č ~� Č ~� � z� � z� Č +  ,VR_NO_BUS       1    ,  O| Č  Y@ Č  Y@ �  O| �  O| Č +  ,VR_NO_BUS       1    ,  �� Č  �@ Č  �@ �  �� �  �� Č +  ,VR_NO_BUS       1    , !�X Č !�@ Č !�@ � !�X � !�X Č +  ,VR_NO_BUS       1    , "�X Č "�@ Č "�@ � "�X � "�X Č +  ,VR_NO_BUS       1    , #�X Č #�@ Č #�@ � #�X � #�X Č +  ,VR_NO_BUS       1    , $�� Č $�@ Č $�@ � $�� � $�� Č +  ,VR_NO_BUS       1    , %� Č %;@ Č %;@ � %� � %� Č +  ,VR_NO_BUS       1    , &1X Č &5@ Č &5@ � &1X � &1X Č +  ,VR_NO_BUS       1    , '+X Č '/@ Č '/@ � '+X � '+X Č +  ,VR_NO_BUS       1    , R( Č m� Č m� � R( � R( Č +  ,VR_NO_BUS       1    , >| Č H@ Č H@ � >| � >| Č +  ,VR_NO_BUS       1    , � Č #  Č #  � � � � Č +  ,VR_NO_BUS       1    ,  Č   Č   �  �  Č +  ,VR_NO_BUS       1    , �� Č �� Č �� � �� � �� Č +  ,VR_NO_BUS       1    , �� Č �� Č �� � �� � �� Č +  ,VR_NO_BUS       1    , Sh Č n� Č n� � Sh � Sh Č +  ,VR_NO_BUS       1    , d� Č h� Č h� � d� � d� Č +  ,VR_NO_BUS       1    , 9� Č C� Č C� � 9� � 9� Č +  ,VR_NO_BUS       1    , 9� Č =� Č =� � 9� � 9� Č +  ,VR_NO_BUS       1    , | Č @ Č @ � | � | Č +  ,VR_NO_BUS       1    , X Č @ Č @ � X � X Č +  ,VR_NO_BUS       1    , �< Č �  Č �  � �< � �< Č +  ,VR_NO_BUS       1    , � Č �  Č �  � � � � Č +  ,VR_NO_BUS       1    , � Č �  Č �  � � � � Č +  ,VR_NO_BUS       1    , .~X �� 0rX �� 0rX �� .~X �� .~X �� +  ,VR_NO_BUS       1    ,  �@ �� Q� �� Q� ��  �@ ��  �@ �� +  ,VR_NO_BUS       1    , �h Č �� Č �� � �h � �h Č +  ,VR_NO_BUS       1    , �� Č �� Č �� � �� � �� Č +  ,VR_NO_BUS       1    , *h Č E� Č E� � *h � *h Č +  ,VR_NO_BUS       1    , � Č  � Č  � � � � � Č +  ,VR_NO_BUS       1    , � Č � Č � � � � � Č +  ,VR_NO_BUS       1    , |( Č �� Č �� � |( � |( Č +  ,VR_NO_BUS       1    , �� Č �� Č �� � �� � �� Č +  ,VR_NO_BUS       1    , b| Č l@ Č l@ � b| � b| Č +  ,VR_NO_BUS       1    , 	bX Č 	f@ Č 	f@ � 	bX � 	bX Č +  ,VR_NO_BUS       1    , 
7< Č 
A  Č 
A  � 
7< � 
7< Č +  ,VR_NO_BUS       1    , 7 Č ;  Č ;  � 7 � 7 Č +  ,VR_NO_BUS       1    , � Č � Č � � � � � Č +  ,VR_NO_BUS       1    , � Č �� Č �� � � � � Č +  ,VR_NO_BUS       1    , "C| �� "M@ �� "M@ �� "C| �� "C| �� +  ,VR_NO_BUS       1    , "�� �� "�@ �� "�@ �� "�� �� "�� �� +  ,VR_NO_BUS       1    , #�< �� #�  �� #�  �� #�< �� #�< �� +  ,VR_NO_BUS       1    , $� �� $"  �� $"  �� $� �� $� �� +  ,VR_NO_BUS       1    , % � �� %  �� %  �� % � �� % � �� +  ,VR_NO_BUS       1    , %�� �� %�@ �� %�@ �� %�� �� %�� �� +  ,VR_NO_BUS       1    , &Xh �� &s� �� &s� �� &Xh �� &Xh �� +  ,VR_NO_BUS       1    , 'i� �� 'm� �� 'm� �� 'i� �� 'i� �� +  ,VR_NO_BUS       1    , (>� �� (H� �� (H� �� (>� �� (>� �� +  ,VR_NO_BUS       1    , )>� �� )B� �� )B� �� )>� �� )>� �� +  ,VR_NO_BUS       1    , *| �� *@ �� *@ �� *| �� *| �� +  ,VR_NO_BUS       1    , *�� �� +@ �� +@ �� *�� �� *�� �� +  ,VR_NO_BUS       1    , ,X �� ,@ �� ,@ �� ,X �� ,X �� +  ,VR_NO_BUS       1    , ,�� �� -@ �� -@ �� ,�� �� ,�� �� +  ,VR_NO_BUS       1    , -l� �� -�@ �� -�@ �� -l� �� -l� �� +  ,VR_NO_BUS       1    , �X �� �@ �� �@ �� �X �� �X �� +  ,VR_NO_BUS       1    , r< �� |  �� |  �� r< �� r< �� +  ,VR_NO_BUS       1    , r �� v  �� v  �� r �� r �� +  ,VR_NO_BUS       1    , l �� p  �� p  �� l �� l �� +  ,VR_NO_BUS       1    , Ѩ �� �  �� �  �� Ѩ �� Ѩ �� +  ,VR_NO_BUS       1    , � �� �  �� �  �� � �� � �� +  ,VR_NO_BUS       1    , � �� �  �� �  �� � �� � �� +  ,VR_NO_BUS       1    , � �� �  �� �  �� � �� � �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �h �� �� �� �� �� �h �� �h �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , z� �� �� �� �� �� z� �� z� �� +  ,VR_NO_BUS       1    , z� �� ~� �� ~� �� z� �� z� �� +  ,VR_NO_BUS       1    ,  t� ��  x� ��  x� ��  t� ��  t� �� +  ,VR_NO_BUS       1    , !n� �� !r� �� !r� �� !n� �� !n� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , 	�� �� 	�� �� 	�� �� 	�� �� 	�� �� +  ,VR_NO_BUS       1    , 
u� �� 
� �� 
� �� 
u� �� 
u� �� +  ,VR_NO_BUS       1    , u� �� y� �� y� �� u� �� u� �� +  ,VR_NO_BUS       1    , 8� �� T@ �� T@ �� 8� �� 8� �� +  ,VR_NO_BUS       1    , JX �� N@ �� N@ �� JX �� JX �� +  ,VR_NO_BUS       1    , DX �� H@ �� H@ �� DX �� DX �� +  ,VR_NO_BUS       1    , �� �� �@ �� �@ �� �� �� �� �� +  ,VR_NO_BUS       1    , �< �� �  �� �  �� �< �� �< �� +  ,VR_NO_BUS       1    , � �� �  �� �  �� � �� � �� +  ,VR_NO_BUS       1    , �� ��   ��   �� �� �� �� �� +  ,VR_NO_BUS       1    ,  ��   ��   ��  ��  �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �@ �� �@ �� �� �� �� �� +  ,VR_NO_BUS       1    , (�( v� (ŀ v� (ŀ � (�( � (�( v� +  ,VR_NO_BUS       1    , )e� v� )�  v� )�  � )e� � )e� v� +  ,VR_NO_BUS       1    , *� v� *@ v� *@ � *� � *� v� +  ,VR_NO_BUS       1    , *~� v� *�@ v� *�@ � *~� � *~� v� +  ,VR_NO_BUS       1    , +�X v� +�@ v� +�@ � +�X � +�X v� +  ,VR_NO_BUS       1    , +�� v� ,@ v� ,@ � +�� � +�� v� +  ,VR_NO_BUS       1    , ,Ш v� ,�  v� ,�  � ,Ш � ,Ш v� +  ,VR_NO_BUS       1    , -� v� 0rX v� 0rX � -� � -� v� +  ,VR_NO_BUS       1    ,  �@ v� Q� v� Q� �  �@ �  �@ v� +  ,VR_NO_BUS       1    , "� �� ,� �� ,� �� "� �� "� �� +  ,VR_NO_BUS       1    , �( �� �� �� �� �� �( �� �( �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , t| �� ~@ �� ~@ �� t| �� t| �� +  ,VR_NO_BUS       1    , �� �� �@ �� �@ �� �� �� �� �� +  ,VR_NO_BUS       1    , �< �� �  �� �  �� �< �� �< �� +  ,VR_NO_BUS       1    , U� v� q@ v� q@ � U� � U� v� +  ,VR_NO_BUS       1    , gX v� k@ v� k@ � gX � gX v� +  ,VR_NO_BUS       1    , aX v� e@ v� e@ � aX � aX v� +  ,VR_NO_BUS       1    , $� v� @  v� @  � $� � $� v� +  ,VR_NO_BUS       1    ,  � v�  � v�  � �  � �  � v� +  ,VR_NO_BUS       1    ,  |h v�  �� v�  �� �  |h �  |h v� +  ,VR_NO_BUS       1    , !�� v� !�� v� !�� � !�� � !�� v� +  ,VR_NO_BUS       1    , "b� v� "l� v� "l� � "b� � "b� v� +  ,VR_NO_BUS       1    , "�( v� "� v� "� � "�( � "�( v� +  ,VR_NO_BUS       1    , #ߘ v� #� v� #� � #ߘ � #ߘ v� +  ,VR_NO_BUS       1    , $٘ v� $݀ v� $݀ � $٘ � $٘ v� +  ,VR_NO_BUS       1    , %?( v� %Z� v� %Z� � %?( � %?( v� +  ,VR_NO_BUS       1    , &9( v� &T� v� &T� � &9( � &9( v� +  ,VR_NO_BUS       1    , 'J� v� 'N� v� 'N� � 'J� � 'J� v� +  ,VR_NO_BUS       1    , '� v� (
  v� (
  � '� � '� v� +  ,VR_NO_BUS       1    , >X v� B@ v� B@ � >X � >X v� +  ,VR_NO_BUS       1    , < v�   v�   � < � < v� +  ,VR_NO_BUS       1    ,  v�   v�   �  �  v� +  ,VR_NO_BUS       1    ,  v�   v�   �  �  v� +  ,VR_NO_BUS       1    , �� v� �� v� �� � �� � �� v� +  ,VR_NO_BUS       1    , �� v� �@ v� �@ � �� � �� v� +  ,VR_NO_BUS       1    , x< v� �  v� �  � x< � x< v� +  ,VR_NO_BUS       1    , x v� |  v� |  � x � x v� +  ,VR_NO_BUS       1    , L� v� V� v� V� � L� � L� v� +  ,VR_NO_BUS       1    , L� v� P� v� P� � L� � L� v� +  ,VR_NO_BUS       1    , !� v� +� v� +� � !� � !� v� +  ,VR_NO_BUS       1    , !� v� %� v� %� � !� � !� v� +  ,VR_NO_BUS       1    , �| v�  @ v�  @ � �| � �| v� +  ,VR_NO_BUS       1    , �X v� �@ v� �@ � �X � �X v� +  ,VR_NO_BUS       1    , �X v� �@ v� �@ � �X � �X v� +  ,VR_NO_BUS       1    , .?� /  0rX /  0rX V .?� V .?� /  +  ,VR_NO_BUS       1    ,  �@ /  Q� /  Q� V  �@ V  �@ /  +  ,VR_NO_BUS       1    , "� v� ,� v� ,� � "� � "� v� +  ,VR_NO_BUS       1    , "� v� &� v� &� � "� � "� v� +  ,VR_NO_BUS       1    , �| v� @ v� @ � �| � �| v� +  ,VR_NO_BUS       1    , �X v� �@ v� �@ � �X � �X v� +  ,VR_NO_BUS       1    , �< v� �  v� �  � �< � �< v� +  ,VR_NO_BUS       1    , � v� �  v� �  � � � � v� +  ,VR_NO_BUS       1    , �� v� �� v� �� � �� � �� v� +  ,VR_NO_BUS       1    , 	�� v� 	�� v� 	�� � 	�� � 	�� v� +  ,VR_NO_BUS       1    , 
�� v� 
�� v� 
�� � 
�� � 
�� v� +  ,VR_NO_BUS       1    , o� v� y� v� y� � o� � o� v� +  ,VR_NO_BUS       1    , o� v� s� v� s� � o� � o� v� +  ,VR_NO_BUS       1    , i� v� m� v� m� � i� � i� v� +  ,VR_NO_BUS       1    , >| v� H@ v� H@ � >| � >| v� +  ,VR_NO_BUS       1    , !�< /  !�  /  !�  V !�< V !�< /  +  ,VR_NO_BUS       1    , "1� /  "M@ /  "M@ V "1� V "1� /  +  ,VR_NO_BUS       1    , #CX /  #G@ /  #G@ V #CX V #CX /  +  ,VR_NO_BUS       1    , #�h /  $� /  $� V #�h V #�h /  +  ,VR_NO_BUS       1    , $�� /  $�  /  $�  V $�� V $�� /  +  ,VR_NO_BUS       1    , %� /  %�  /  %�  V %� V %� /  +  ,VR_NO_BUS       1    , &i� /  &s� /  &s� V &i� V &i� /  +  ,VR_NO_BUS       1    , 'i� /  'm� /  'm� V 'i� V 'i� /  +  ,VR_NO_BUS       1    , '� /  (
  /  (
  V '� V '� /  +  ,VR_NO_BUS       1    , )  /  )  /  )  V )  V )  /  +  ,VR_NO_BUS       1    , )� /  )�  /  )�  V )� V )� /  +  ,VR_NO_BUS       1    , *~� /  *�@ /  *�@ V *~� V *~� /  +  ,VR_NO_BUS       1    , +:h /  +U� /  +U� V +:h V +:h /  +  ,VR_NO_BUS       1    , ,K� /  ,O� /  ,O� V ,K� V ,K� /  +  ,VR_NO_BUS       1    , - � /  -I� /  -I� V - � V - � /  +  ,VR_NO_BUS       1    , �< /  �  /  �  V �< V �< /  +  ,VR_NO_BUS       1    , Z� /  v  /  v  V Z� V Z� /  +  ,VR_NO_BUS       1    , l /  p  /  p  V l V l /  +  ,VR_NO_BUS       1    , @� /  J� /  J� V @� V @� /  +  ,VR_NO_BUS       1    , �h /  �� /  �� V �h V �h /  +  ,VR_NO_BUS       1    , �� /  �� /  �� V �� V �� /  +  ,VR_NO_BUS       1    , #h /  >� /  >� V #h V #h /  +  ,VR_NO_BUS       1    , �( /  � /  � V �( V �( /  +  ,VR_NO_BUS       1    , � /  � /  � V � V � /  +  ,VR_NO_BUS       1    , �h /  �� /  �� V �h V �h /  +  ,VR_NO_BUS       1    , O� /  k@ /  k@ V O� V O� /  +  ,VR_NO_BUS       1    , aX /  e@ /  e@ V aX V aX /  +  ,VR_NO_BUS       1    , 6< /  @  /  @  V 6< V 6< /  +  ,VR_NO_BUS       1    , �� /  �@ /  �@ V �� V �� /  +  ,VR_NO_BUS       1    ,  �X /   �@ /   �@ V  �X V  �X /  +  ,VR_NO_BUS       1    , 	�� /  	�  /  	�  V 	�� V 	�� /  +  ,VR_NO_BUS       1    , 
� /  
�  /  
�  V 
� V 
� /  +  ,VR_NO_BUS       1    , � /  ;  /  ;  V � V � /  +  ,VR_NO_BUS       1    , � /  � /  � V � V � /  +  ,VR_NO_BUS       1    , � /  �� /  �� V � V � /  +  ,VR_NO_BUS       1    , �| /  �@ /  �@ V �| V �| /  +  ,VR_NO_BUS       1    , ,� /  H@ /  H@ V ,� V ,� /  +  ,VR_NO_BUS       1    , �� /  �@ /  �@ V �� V �� /  +  ,VR_NO_BUS       1    , �< /  �  /  �  V �< V �< /  +  ,VR_NO_BUS       1    , p� /  z� /  z� V p� V p� /  +  ,VR_NO_BUS       1    , p� /  t� /  t� V p� V p� /  +  ,VR_NO_BUS       1    , E� /  O� /  O� V E� V E� /  +  ,VR_NO_BUS       1    , E� /  I� /  I� V E� V E� /  +  ,VR_NO_BUS       1    , | /  $@ /  $@ V | V | /  +  ,VR_NO_BUS       1    , X /  @ /  @ V X V X /  +  ,VR_NO_BUS       1    , +Q� 
ɸ +�@ 
ɸ +�@ 
�� +Q� 
�� +Q� 
ɸ +  ,VR_NO_BUS       1    , ,4h 
ɸ ,O� 
ɸ ,O� 
�� ,4h 
�� ,4h 
ɸ +  ,VR_NO_BUS       1    , ,Ш 
ɸ ,�  
ɸ ,�  
�� ,Ш 
�� ,Ш 
ɸ +  ,VR_NO_BUS       1    , -� 
ɸ -�  
ɸ -�  
�� -� 
�� -� 
ɸ +  ,VR_NO_BUS       1    , .f� 
ɸ 0rX 
ɸ 0rX 
�� .f� 
�� .f� 
ɸ +  ,VR_NO_BUS       1    ,  �@ 
ɸ Q� 
ɸ Q� 
��  �@ 
��  �@ 
ɸ +  ,VR_NO_BUS       1    , Ҩ /  �  /  �  V Ҩ V Ҩ /  +  ,VR_NO_BUS       1    , � /  �  /  �  V � V � /  +  ,VR_NO_BUS       1    , �h /  �� /  �� V �h V �h /  +  ,VR_NO_BUS       1    , $h /  ?� /  ?� V $h V $h /  +  ,VR_NO_BUS       1    , �( /  � /  � V �( V �( /  +  ,VR_NO_BUS       1    , � /  � /  � V � V � /  +  ,VR_NO_BUS       1    , �� /  �  /  �  V �� V �� /  +  ,VR_NO_BUS       1    , P� /  l@ /  l@ V P� V P� /  +  ,VR_NO_BUS       1    , 	=< /  	G  /  	G  V 	=< V 	=< /  +  ,VR_NO_BUS       1    , aX 
ɸ e@ 
ɸ e@ 
�� aX 
�� aX 
ɸ +  ,VR_NO_BUS       1    , [X 
ɸ _@ 
ɸ _@ 
�� [X 
�� [X 
ɸ +  ,VR_NO_BUS       1    , �h 
ɸ  � 
ɸ  � 
�� �h 
�� �h 
ɸ +  ,VR_NO_BUS       1    ,  �� 
ɸ  �@ 
ɸ  �@ 
��  �� 
��  �� 
ɸ +  ,VR_NO_BUS       1    , !�X 
ɸ !�@ 
ɸ !�@ 
�� !�X 
�� !�X 
ɸ +  ,VR_NO_BUS       1    , "�� 
ɸ "�@ 
ɸ "�@ 
�� "�� 
�� "�� 
ɸ +  ,VR_NO_BUS       1    , #+� 
ɸ #G@ 
ɸ #G@ 
�� #+� 
�� #+� 
ɸ +  ,VR_NO_BUS       1    , $=X 
ɸ $A@ 
ɸ $A@ 
�� $=X 
�� $=X 
ɸ +  ,VR_NO_BUS       1    , $�( 
ɸ $݀ 
ɸ $݀ 
�� $�( 
�� $�( 
ɸ +  ,VR_NO_BUS       1    , %�| 
ɸ %�@ 
ɸ %�@ 
�� %�| 
�� %�| 
ɸ +  ,VR_NO_BUS       1    , &�< 
ɸ &�  
ɸ &�  
�� &�< 
�� &�< 
ɸ +  ,VR_NO_BUS       1    , '� 
ɸ '�  
ɸ '�  
�� '� 
�� '� 
ɸ +  ,VR_NO_BUS       1    , (� 
ɸ (�  
ɸ (�  
�� (� 
�� (� 
ɸ +  ,VR_NO_BUS       1    , )W� 
ɸ )a� 
ɸ )a� 
�� )W� 
�� )W� 
ɸ +  ,VR_NO_BUS       1    , *W� 
ɸ *[� 
ɸ *[� 
�� *W� 
�� *W� 
ɸ +  ,VR_NO_BUS       1    , �\ 
ɸ �� 
ɸ �� 
�� �\ 
�� �\ 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �@ 
ɸ �@ 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �@ 
ɸ �@ 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , �( 
ɸ ƀ 
ɸ ƀ 
�� �( 
�� �( 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �� 
ɸ �� 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , �| 
ɸ �@ 
ɸ �@ 
�� �| 
�� �| 
ɸ +  ,VR_NO_BUS       1    , l< 
ɸ v  
ɸ v  
�� l< 
�� l< 
ɸ +  ,VR_NO_BUS       1    , ר 
ɸ �  
ɸ �  
�� ר 
�� ר 
ɸ +  ,VR_NO_BUS       1    , � 
ɸ �  
ɸ �  
�� � 
�� � 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �� 
ɸ �� 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �� 
ɸ �� 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �� 
ɸ �� 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �� 
ɸ �� 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �� 
ɸ �� 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , a| 
ɸ k@ 
ɸ k@ 
�� a| 
�� a| 
ɸ +  ,VR_NO_BUS       1    , �( 
ɸ �� 
ɸ �� 
�� �( 
�� �( 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ �� 
ɸ �� 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , h 
ɸ 9� 
ɸ 9� 
�� h 
�� h 
ɸ +  ,VR_NO_BUS       1    , 
� 
ɸ � 
ɸ � 
�� 
� 
�� 
� 
ɸ +  ,VR_NO_BUS       1    , 
� 
ɸ � 
ɸ � 
�� 
� 
�� 
� 
ɸ +  ,VR_NO_BUS       1    , �h 
ɸ �� 
ɸ �� 
�� �h 
�� �h 
ɸ +  ,VR_NO_BUS       1    , 	�\ 
ɸ 	�� 
ɸ 	�� 
�� 	�\ 
�� 	�\ 
ɸ +  ,VR_NO_BUS       1    , 
�\ 
ɸ 
�� 
ɸ 
�� 
�� 
�\ 
�� 
�\ 
ɸ +  ,VR_NO_BUS       1    , o� 
ɸ y� 
ɸ y� 
�� o� 
�� o� 
ɸ +  ,VR_NO_BUS       1    , �( 
ɸ �� 
ɸ �� 
�� �( 
�� �( 
ɸ +  ,VR_NO_BUS       1    , �| 
ɸ �@ 
ɸ �@ 
�� �| 
�� �| 
ɸ +  ,VR_NO_BUS       1    , T 
ɸ m� 
ɸ m� 
�� T 
�� T 
ɸ +  ,VR_NO_BUS       1    , �\ 
ɸ 	� 
ɸ 	� 
�� �\ 
�� �\ 
ɸ +  ,VR_NO_BUS       1    , ڼ 
ɸ � 
ɸ � 
�� ڼ 
�� ڼ 
ɸ +  ,VR_NO_BUS       1    , �h 
ɸ �� 
ɸ �� 
�� �h 
�� �h 
ɸ +  ,VR_NO_BUS       1    , $�X � $�@ � $�@ � $�X � $�X � +  ,VR_NO_BUS       1    , %}� � %�  � %�  � %}� � %}� � +  ,VR_NO_BUS       1    , &9( � &T� � &T� � &9( � &9( � +  ,VR_NO_BUS       1    , &�( � &р � &р � &�( � &�( � +  ,VR_NO_BUS       1    , 'ǘ � 'ˀ � 'ˀ � 'ǘ � 'ǘ � +  ,VR_NO_BUS       1    , (�| � (�@ � (�@ � (�| � (�| � +  ,VR_NO_BUS       1    , )w< � )�  � )�  � )w< � )w< � +  ,VR_NO_BUS       1    , *w � *{  � *{  � *w � *w � +  ,VR_NO_BUS       1    , +q � +u  � +u  � +q � +q � +  ,VR_NO_BUS       1    , ,k � ,o  � ,o  � ,k � ,k � +  ,VR_NO_BUS       1    , -e � -i  � -i  � -e � -e � +  ,VR_NO_BUS       1    , .9� � 0rX � 0rX � .9� � .9� � +  ,VR_NO_BUS       1    ,  �@ � Q� � Q� �  �@ �  �@ � +  ,VR_NO_BUS       1    , G� 
ɸ K� 
ɸ K� 
�� G� 
�� G� 
ɸ +  ,VR_NO_BUS       1    , �� 
ɸ @ 
ɸ @ 
�� �� 
�� �� 
ɸ +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , m| � w@ � w@ � m| � m| � +  ,VR_NO_BUS       1    , H< � R  � R  � H< � H< � +  ,VR_NO_BUS       1    , "� � ,� � ,� � "� � "� � +  ,VR_NO_BUS       1    , "� � &� � &� � "� � "� � +  ,VR_NO_BUS       1    , �� � �@ � �@ � �� � �� � +  ,VR_NO_BUS       1    , �h � �� � �� � �h � �h � +  ,VR_NO_BUS       1    ,  n� �  x� �  x� �  n� �  n� � +  ,VR_NO_BUS       1    , !n� � !r� � !r� � !n� � !n� � +  ,VR_NO_BUS       1    , "C| � "M@ � "M@ � "C| � "C| � +  ,VR_NO_BUS       1    , #CX � #G@ � #G@ � #CX � #CX � +  ,VR_NO_BUS       1    , #�� � #�@ � #�@ � #�� � #�� � +  ,VR_NO_BUS       1    , �� � �@ � �@ � �� � �� � +  ,VR_NO_BUS       1    , 2� � N@ � N@ � 2� � 2� � +  ,VR_NO_BUS       1    , �� � �@ � �@ � �� � �� � +  ,VR_NO_BUS       1    , �( � � � � � �( � �( � +  ,VR_NO_BUS       1    , �� � �@ � �@ � �� � �� � +  ,VR_NO_BUS       1    ,  � � <@ � <@ �  � �  � � +  ,VR_NO_BUS       1    , < �   �   � < � < � +  ,VR_NO_BUS       1    , x� � �  � �  � x� � x� � +  ,VR_NO_BUS       1    , �� �   �   � �� � �� � +  ,VR_NO_BUS       1    , � � ̀ � ̀ � � � � � +  ,VR_NO_BUS       1    , �| � �@ � �@ � �| � �| � +  ,VR_NO_BUS       1    , � � $@ � $@ � � � � � +  ,VR_NO_BUS       1    , � � @ � @ � � � � � +  ,VR_NO_BUS       1    , �< � �  � �  � �< � �< � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , ,�� tX ,�� tX ,�� �h ,�� �h ,�� tX +  ,VR_NO_BUS       1    , -~| tX -�@ tX -�@ �h -~| �h -~| tX +  ,VR_NO_BUS       1    , .~X tX 0rX tX 0rX �h .~X �h .~X tX +  ,VR_NO_BUS       1    ,  �@ tX Q� tX Q� �h  �@ �h  �@ tX +  ,VR_NO_BUS       1    , Ҩ � �  � �  � Ҩ � Ҩ � +  ,VR_NO_BUS       1    , � � �  � �  � � � � � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , b| � l@ � l@ � b| � b| � +  ,VR_NO_BUS       1    , 	=< � 	G  � 	G  � 	=< � 	=< � +  ,VR_NO_BUS       1    , 
D� � 
`@ � 
`@ � 
D� � 
D� � +  ,VR_NO_BUS       1    , 
�� � 
�@ � 
�@ � 
�� � 
�� � +  ,VR_NO_BUS       1    , �( � �� � �� � �( � �( � +  ,VR_NO_BUS       1    , � tX  � tX  � �h � �h � tX +  ,VR_NO_BUS       1    ,  � tX  � tX  � �h  � �h  � tX +  ,VR_NO_BUS       1    ,  � tX  �� tX  �� �h  � �h  � tX +  ,VR_NO_BUS       1    , !� tX !� tX !� �h !� �h !� tX +  ,VR_NO_BUS       1    , "�| tX "�@ tX "�@ �h "�| �h "�| tX +  ,VR_NO_BUS       1    , #�X tX #�@ tX #�@ �h #�X �h #�X tX +  ,VR_NO_BUS       1    , $�X tX $�@ tX $�@ �h $�X �h $�X tX +  ,VR_NO_BUS       1    , %�X tX %�@ tX %�@ �h %�X �h %�X tX +  ,VR_NO_BUS       1    , &w� tX &�  tX &�  �h &w� �h &w� tX +  ,VR_NO_BUS       1    , '� tX '�  tX '�  �h '� �h '� tX +  ,VR_NO_BUS       1    , (]� tX (g� tX (g� �h (]� �h (]� tX +  ,VR_NO_BUS       1    , )]� tX )a� tX )a� �h )]� �h )]� tX +  ,VR_NO_BUS       1    , )� tX )�  tX )�  �h )� �h )� tX +  ,VR_NO_BUS       1    , *�� tX *�� tX *�� �h *�� �h *�� tX +  ,VR_NO_BUS       1    , +�� tX +�� tX +�� �h +�� �h +�� tX +  ,VR_NO_BUS       1    , 4( tX O� tX O� �h 4( �h 4( tX +  ,VR_NO_BUS       1    , � tX *@ tX *@ �h � �h � tX +  ,VR_NO_BUS       1    , (( tX C� tX C� �h (( �h (( tX +  ,VR_NO_BUS       1    , �( tX �� tX �� �h �( �h �( tX +  ,VR_NO_BUS       1    , �h tX �� tX �� �h �h �h �h tX +  ,VR_NO_BUS       1    , �( tX �� tX �� �h �( �h �( tX +  ,VR_NO_BUS       1    , �h tX �� tX �� �h �h �h �h tX +  ,VR_NO_BUS       1    , /h tX J� tX J� �h /h �h /h tX +  ,VR_NO_BUS       1    , � tX %� tX %� �h � �h � tX +  ,VR_NO_BUS       1    , �| tX  @ tX  @ �h �| �h �| tX +  ,VR_NO_BUS       1    , �< tX �  tX �  �h �< �h �< tX +  ,VR_NO_BUS       1    , � tX �  tX �  �h � �h � tX +  ,VR_NO_BUS       1    , � tX �  tX �  �h � �h � tX +  ,VR_NO_BUS       1    , �� tX �� tX �� �h �� �h �� tX +  ,VR_NO_BUS       1    , *� tX F  tX F  �h *� �h *� tX +  ,VR_NO_BUS       1    , �� tX �  tX �  �h �� �h �� tX +  ,VR_NO_BUS       1    , �� tX �� tX �� �h �� �h �� tX +  ,VR_NO_BUS       1    , 	�� tX 	�� tX 	�� �h 	�� �h 	�� tX +  ,VR_NO_BUS       1    , 
�� tX 
�  tX 
�  �h 
�� �h 
�� tX +  ,VR_NO_BUS       1    , ^( tX y� tX y� �h ^( �h ^( tX +  ,VR_NO_BUS       1    , �( tX �� tX �� �h �( �h �( tX +  ,VR_NO_BUS       1    , �| tX �@ tX �@ �h �| �h �| tX +  ,VR_NO_BUS       1    , �< tX �  tX �  �h �< �h �< tX +  ,VR_NO_BUS       1    , � tX �  tX �  �h � �h � tX +  ,VR_NO_BUS       1    , � tX #  tX #  �h � �h � tX +  ,VR_NO_BUS       1    , �� tX �@ tX �@ �h �� �h �� tX +  ,VR_NO_BUS       1    ,  � tX <@ tX <@ �h  � �h  � tX +  ,VR_NO_BUS       1    , �( tX ؀ tX ؀ �h �( �h �( tX +  ,VR_NO_BUS       1    , :( tX U� tX U� �h :( �h :( tX +  ,VR_NO_BUS       1    , �( tX Ҁ tX Ҁ �h �( �h �( tX +  ,VR_NO_BUS       1    , (%X l� ()@ l� ()@ �� (%X �� (%X l� +  ,VR_NO_BUS       1    , )X l� )#@ l� )#@ �� )X �� )X l� +  ,VR_NO_BUS       1    , )�( l� )�� l� )�� �� )�( �� )�( l� +  ,VR_NO_BUS       1    , *_� l� *{  l� *{  �� *_� �� *_� l� +  ,VR_NO_BUS       1    , *�� l� +@ l� +@ �� *�� �� *�� l� +  ,VR_NO_BUS       1    , +�h l� +�� l� +�� �� +�h �� +�h l� +  ,VR_NO_BUS       1    , ,r� l� ,�@ l� ,�@ �� ,r� �� ,r� l� +  ,VR_NO_BUS       1    , -.h l� 0rX l� 0rX �� -.h �� -.h l� +  ,VR_NO_BUS       1    ,  �@ l� Q� l� Q� ��  �@ ��  �@ l� +  ,VR_NO_BUS       1    , Ҩ tX �  tX �  �h Ҩ �h Ҩ tX +  ,VR_NO_BUS       1    , �� tX �� tX �� �h �� �h �� tX +  ,VR_NO_BUS       1    , �� tX �� tX �� �h �� �h �� tX +  ,VR_NO_BUS       1    , �� tX �� tX �� �h �� �h �� tX +  ,VR_NO_BUS       1    , n| tX x@ tX x@ �h n| �h n| tX +  ,VR_NO_BUS       1    , I< tX S  tX S  �h I< �h I< tX +  ,VR_NO_BUS       1    , �h l� �� l� �� �� �h �� �h l� +  ,VR_NO_BUS       1    , 6� l� R  l� R  �� 6� �� 6� l� +  ,VR_NO_BUS       1    , "� l� ,� l� ,� �� "� �� "� l� +  ,VR_NO_BUS       1    , "� l� &� l� &� �� "� �� "� l� +  ,VR_NO_BUS       1    , � l�  � l�  � �� � �� � l� +  ,VR_NO_BUS       1    , � l� �� l� �� �� � �� � l� +  ,VR_NO_BUS       1    ,  � l�  �� l�  �� ��  � ��  � l� +  ,VR_NO_BUS       1    , !� l� !� l� !� �� !� �� !� l� +  ,VR_NO_BUS       1    , "�| l� "�@ l� "�@ �� "�| �� "�| l� +  ,VR_NO_BUS       1    , #�< l� #�  l� #�  �� #�< �� #�< l� +  ,VR_NO_BUS       1    , $%� l� $A@ l� $A@ �� $%� �� $%� l� +  ,VR_NO_BUS       1    , $�� l� $�@ l� $�@ �� $�� �� $�� l� +  ,VR_NO_BUS       1    , %�X l� %�@ l� %�@ �� %�X �� %�X l� +  ,VR_NO_BUS       1    , &9( l� &T� l� &T� �� &9( �� &9( l� +  ,VR_NO_BUS       1    , '%| l� '/@ l� '/@ �� '%| �� '%| l� +  ,VR_NO_BUS       1    , � l� �  l� �  �� � �� � l� +  ,VR_NO_BUS       1    , p� l� z� l� z� �� p� �� p� l� +  ,VR_NO_BUS       1    , � l� 6@ l� 6@ �� � �� � l� +  ,VR_NO_BUS       1    , �� l� �@ l� �@ �� �� �� �� l� +  ,VR_NO_BUS       1    , �X l� �@ l� �@ �� �X �� �X l� +  ,VR_NO_BUS       1    , ~< l� �  l� �  �� ~< �� ~< l� +  ,VR_NO_BUS       1    , ~ l� �  l� �  �� ~ �� ~ l� +  ,VR_NO_BUS       1    , R� l� \� l� \� �� R� �� R� l� +  ,VR_NO_BUS       1    , R� l� V� l� V� �� R� �� R� l� +  ,VR_NO_BUS       1    , L� l� P� l� P� �� L� �� L� l� +  ,VR_NO_BUS       1    , �h l� �� l� �� �� �h �� �h l� +  ,VR_NO_BUS       1    , �� l� �� l� �� �� �� �� �� l� +  ,VR_NO_BUS       1    , �� l� �� l� �� �� �� �� �� l� +  ,VR_NO_BUS       1    , B� l� ^  l� ^  �� B� �� B� l� +  ,VR_NO_BUS       1    , .� l� 8� l� 8� �� .� �� .� l� +  ,VR_NO_BUS       1    , G� l� K� l� K� �� G� �� G� l� +  ,VR_NO_BUS       1    , A� l� E� l� E� �� A� �� A� l� +  ,VR_NO_BUS       1    , ( l�  � l�  � �� ( �� ( l� +  ,VR_NO_BUS       1    , �( l� �� l� �� �� �( �� �( l� +  ,VR_NO_BUS       1    , n| l� x@ l� x@ �� n| �� n| l� +  ,VR_NO_BUS       1    , nX l� r@ l� r@ �� nX �� nX l� +  ,VR_NO_BUS       1    , C< l� M  l� M  �� C< �� C< l� +  ,VR_NO_BUS       1    , 	� l� 	'� l� 	'� �� 	� �� 	� l� +  ,VR_NO_BUS       1    , 
� l� 
!� l� 
!� �� 
� �� 
� l� +  ,VR_NO_BUS       1    , 
�h l� 
�� l� 
�� �� 
�h �� 
�h l� +  ,VR_NO_BUS       1    ,  h l� � l� � ��  h ��  h l� +  ,VR_NO_BUS       1    , � l� �� l� �� �� � �� � l� +  ,VR_NO_BUS       1    , � l� �� l� �� �� � �� � l� +  ,VR_NO_BUS       1    , �| l� �@ l� �@ �� �| �� �| l� +  ,VR_NO_BUS       1    , �< l� �  l� �  �� �< �� �< l� +  ,VR_NO_BUS       1    , !*< "� !4  "� !4  I� !*< I� !*< "� +  ,VR_NO_BUS       1    , "* "� ".  "� ".  I� "* I� "* "� +  ,VR_NO_BUS       1    , #$ "� #(  "� #(  I� #$ I� #$ "� +  ,VR_NO_BUS       1    , #�h "� $� "� $� I� #�h I� #�h "� +  ,VR_NO_BUS       1    , $dh "� $� "� $� I� $dh I� $dh "� +  ,VR_NO_BUS       1    , %u� "� %y� "� %y� I� %u� I� %u� "� +  ,VR_NO_BUS       1    , &� "� &5@ "� &5@ I� &� I� &� "� +  ,VR_NO_BUS       1    , '+X "� '/@ "� '/@ I� '+X I� '+X "� +  ,VR_NO_BUS       1    , ( < "� (
  "� (
  I� ( < I� ( < "� +  ,VR_NO_BUS       1    , )  "� )  "� )  I� )  I� )  "� +  ,VR_NO_BUS       1    , )�� "� )�@ "� )�@ I� )�� I� )�� "� +  ,VR_NO_BUS       1    , *@h "� *[� "� *[� I� *@h I� *@h "� +  ,VR_NO_BUS       1    , *�� "� +@ "� +@ I� *�� I� *�� "� +  ,VR_NO_BUS       1    , ,X "� 0rX "� 0rX I� ,X I� ,X "� +  ,VR_NO_BUS       1    ,  �@ "� Q� "� Q� I�  �@ I�  �@ "� +  ,VR_NO_BUS       1    , X� "� b� "� b� I� X� I� X� "� +  ,VR_NO_BUS       1    , 3� "� =� "� =� I� 3� I� 3� "� +  ,VR_NO_BUS       1    , �( "� �� "� �� I� �( I� �( "� +  ,VR_NO_BUS       1    , �� "� �� "� �� I� �� I� �� "� +  ,VR_NO_BUS       1    , �� "� �� "� �� I� �� I� �� "� +  ,VR_NO_BUS       1    , /h "� J� "� J� I� /h I� /h "� +  ,VR_NO_BUS       1    , � "� %� "� %� I� � I� � "� +  ,VR_NO_BUS       1    , �| "�  @ "�  @ I� �| I� �| "� +  ,VR_NO_BUS       1    , �< "� �  "� �  I� �< I� �< "� +  ,VR_NO_BUS       1    , � "� �  "� �  I� � I� � "� +  ,VR_NO_BUS       1    , �� "� �� "� �� I� �� I� �� "� +  ,VR_NO_BUS       1    , �� "� �� "� �� I� �� I� �� "� +  ,VR_NO_BUS       1    , z� "� �� "� �� I� z� I� z� "� +  ,VR_NO_BUS       1    , U| "� _@ "� _@ I� U| I� U| "� +  ,VR_NO_BUS       1    ,  UX "�  Y@ "�  Y@ I�  UX I�  UX "� +  ,VR_NO_BUS       1    , �� "� �@ "� �@ I� �� I� �� "� +  ,VR_NO_BUS       1    , �X "� �@ "� �@ I� �X I� �X "� +  ,VR_NO_BUS       1    , 	�< "� 	�  "� 	�  I� 	�< I� 	�< "� +  ,VR_NO_BUS       1    , 
� "� 
�  "� 
�  I� 
� I� 
� "� +  ,VR_NO_BUS       1    , �� "� �� "� �� I� �� I� �� "� +  ,VR_NO_BUS       1    , �h "� � "� � I� �h I� �h "� +  ,VR_NO_BUS       1    , � "� � "� � I� � I� � "� +  ,VR_NO_BUS       1    , � "� 	� "� 	� I� � I� � "� +  ,VR_NO_BUS       1    , kh "� �� "� �� I� kh I� kh "� +  ,VR_NO_BUS       1    , W� "� a� "� a� I� W� I� W� "� +  ,VR_NO_BUS       1    , 2| "� <@ "� <@ I� 2| I� 2| "� +  ,VR_NO_BUS       1    , 2X "� 6@ "� 6@ I� 2X I� 2X "� +  ,VR_NO_BUS       1    , < "�   "�   I� < I� < "� +  ,VR_NO_BUS       1    , r� "� �  "� �  I� r� I� r� "� +  ,VR_NO_BUS       1    , � "� �  "� �  I� � I� � "� +  ,VR_NO_BUS       1    , %u�  X %y�  X %y�  Bh %u�  Bh %u�  X +  ,VR_NO_BUS       1    , &o�  X &s�  X &s�  Bh &o�  Bh &o�  X +  ,VR_NO_BUS       1    , &��  X '   X '   Bh &��  Bh &��  X +  ,VR_NO_BUS       1    , '��  X '��  X '��  Bh '��  Bh '��  X +  ,VR_NO_BUS       1    , (��  X (ŀ  X (ŀ  Bh (��  Bh (��  X +  ,VR_NO_BUS       1    , )��  X )��  X )��  Bh )��  Bh )��  X +  ,VR_NO_BUS       1    , *_�  X *{   X *{   Bh *_�  Bh *_�  X +  ,VR_NO_BUS       1    , +(  X 0rX  X 0rX  Bh +(  Bh +(  X +  ,VR_NO_BUS       1    ,  �@  X Q�  X Q�  Bh  �@  Bh  �@  X +  ,VR_NO_BUS       1    , G� "� K� "� K� I� G� I� G� "� +  ,VR_NO_BUS       1    , ( "� &� "� &� I� ( I� ( "� +  ,VR_NO_BUS       1    , �( "� �� "� �� I� �( I� �( "� +  ,VR_NO_BUS       1    , �� "� �� "� �� I� �� I� �� "� +  ,VR_NO_BUS       1    , n| "� x@ "� x@ I� n| I� n| "� +  ,VR_NO_BUS       1    , nX "� r@ "� r@ I� nX I� nX "� +  ,VR_NO_BUS       1    , ��  X ��  X ��  Bh ��  Bh ��  X +  ,VR_NO_BUS       1    , ��  X ��  X ��  Bh ��  Bh ��  X +  ,VR_NO_BUS       1    , ��  X ��  X ��  Bh ��  Bh ��  X +  ,VR_NO_BUS       1    , s|  X }@  X }@  Bh s|  Bh s|  X +  ,VR_NO_BUS       1    , sX  X w@  X w@  Bh sX  Bh sX  X +  ,VR_NO_BUS       1    , H<  X R   X R   Bh H<  Bh H<  X +  ,VR_NO_BUS       1    , "�  X ,�  X ,�  Bh "�  Bh "�  X +  ,VR_NO_BUS       1    , ��  X �  X �  Bh ��  Bh ��  X +  ,VR_NO_BUS       1    , ��  X �  X �  Bh ��  Bh ��  X +  ,VR_NO_BUS       1    , ��  X ��  X ��  Bh ��  Bh ��  X +  ,VR_NO_BUS       1    ,  �|  X  �@  X  �@  Bh  �|  Bh  �|  X +  ,VR_NO_BUS       1    , !�X  X !�@  X !�@  Bh !�X  Bh !�X  X +  ,VR_NO_BUS       1    , "�<  X "�   X "�   Bh "�<  Bh "�<  X +  ,VR_NO_BUS       1    , #�  X #�   X #�   Bh #�  Bh #�  X +  ,VR_NO_BUS       1    , $u�  X $�  X $�  Bh $u�  Bh $u�  X +  ,VR_NO_BUS       1    , 
�  X 
!�  X 
!�  Bh 
�  Bh 
�  X +  ,VR_NO_BUS       1    , �  X �  X �  Bh �  Bh �  X +  ,VR_NO_BUS       1    , �(  X ��  X ��  Bh �(  Bh �(  X +  ,VR_NO_BUS       1    , �  X ��  X ��  Bh �  Bh �  X +  ,VR_NO_BUS       1    , �  X �  X �  Bh �  Bh �  X +  ,VR_NO_BUS       1    , �|  X �@  X �@  Bh �|  Bh �|  X +  ,VR_NO_BUS       1    , �<  X �   X �   Bh �<  Bh �<  X +  ,VR_NO_BUS       1    , �  X �   X �   Bh �  Bh �  X +  ,VR_NO_BUS       1    , j�  X t�  X t�  Bh j�  Bh j�  X +  ,VR_NO_BUS       1    , E�  X O�  X O�  Bh E�  Bh E�  X +  ,VR_NO_BUS       1    , E�  X I�  X I�  Bh E�  Bh E�  X +  ,VR_NO_BUS       1    , |  X $@  X $@  Bh |  Bh |  X +  ,VR_NO_BUS       1    , X  X @  X @  Bh X  Bh X  X +  ,VR_NO_BUS       1    , �<  X �   X �   Bh �<  Bh �<  X +  ,VR_NO_BUS       1    , ��  X ��  X ��  Bh ��  Bh ��  X +  ,VR_NO_BUS       1    , #< &�� #(  &�� #(  &�� #< &�� #< &�� +  ,VR_NO_BUS       1    , %�� &�� &  &�� &  &�� %�� &�� %�� &�� +  ,VR_NO_BUS       1    , (� &�� )#@ &�� )#@ &�� (� &�� (� &�� +  ,VR_NO_BUS       1    , �� �� �$ �� �$ �� �� �� �� ��      1    , ! Ӝ #�d Ӝ #�d �T ! �T ! Ӝ      1    , v� � �� � �� x v� x v� �      1    , G�  X K�  X K�  Bh G�  Bh G�  X +  ,VR_NO_BUS       1    , �h  X ��  X ��  Bh �h  Bh �h  X +  ,VR_NO_BUS       1    , �(  X ��  X ��  Bh �(  Bh �(  X +  ,VR_NO_BUS       1    , (  X  �  X  �  Bh (  Bh (  X +  ,VR_NO_BUS       1    , �  X �  X �  Bh �  Bh �  X +  ,VR_NO_BUS       1    , �|  X �@  X �@  Bh �|  Bh �|  X +  ,VR_NO_BUS       1    , �X  X �@  X �@  Bh �X  Bh �X  X +  ,VR_NO_BUS       1    , ��  X �   X �   Bh ��  Bh ��  X +  ,VR_NO_BUS       1    , 	+�  X 	G   X 	G   Bh 	+�  Bh 	+�  X +  ,VR_NO_BUS       1    , X &�� @ &�� @ &�� X &�� X &�� +  ,VR_NO_BUS       1    , �< &�� �  &�� �  &�� �< &�� �< &�� +  ,VR_NO_BUS       1    , � &�� �  &�� �  &�� � &�� � &�� +  ,VR_NO_BUS       1    , � &�� �  &�� �  &�� � &�� � &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , [| &�� e@ &�� e@ &�� [| &�� [| &�� +  ,VR_NO_BUS       1    , [X &�� _@ &�� _@ &�� [X &�� [X &�� +  ,VR_NO_BUS       1    ,  UX &��  Y@ &��  Y@ &��  UX &��  UX &�� +  ,VR_NO_BUS       1    ,  �� &��  �@ &��  �@ &��  �� &��  �� &�� +  ,VR_NO_BUS       1    , !�X &�� !�@ &�� !�@ &�� !�X &�� !�X &�� +  ,VR_NO_BUS       1    , "1� &�� "M@ &�� "M@ &�� "1� &�� "1� &�� +  ,VR_NO_BUS       1    , 	h &�� 	'� &�� 	'� &�� 	h &�� 	h &�� +  ,VR_NO_BUS       1    , 
� &�� 
!� &�� 
!� &�� 
� &�� 
� &�� +  ,VR_NO_BUS       1    , 
�� &�� 
�  &�� 
�  &�� 
�� &�� 
�� &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , ,� &�� H@ &�� H@ &�� ,� &�� ,� &�� +  ,VR_NO_BUS       1    , �h &�� � &�� � &�� �h &�� �h &�� +  ,VR_NO_BUS       1    , Լ &�� ހ &�� ހ &�� Լ &�� Լ &�� +  ,VR_NO_BUS       1    , Ԙ &�� ؀ &�� ؀ &�� Ԙ &�� Ԙ &�� +  ,VR_NO_BUS       1    , :( &�� U� &�� U� &�� :( &�� :( &�� +  ,VR_NO_BUS       1    , K� &�� O� &�� O� &�� K� &�� K� &�� +  ,VR_NO_BUS       1    ,  | &�� *@ &�� *@ &��  | &��  | &�� +  ,VR_NO_BUS       1    ,  X &�� $@ &�� $@ &��  X &��  X &�� +  ,VR_NO_BUS       1    , X &�� @ &�� @ &�� X &�� X &�� +  ,VR_NO_BUS       1    , &J� $�L &T� $�L &T� $�\ &J� $�\ &J� $�L +  ,VR_NO_BUS       1    , 'J� $�L 'N� $�L 'N� $�\ 'J� $�\ 'J� $�L +  ,VR_NO_BUS       1    , *!( $�L *<� $�L *<� $�\ *!( $�\ *!( $�L +  ,VR_NO_BUS       1    , -( $�L -*� $�L -*� $�\ -( $�\ -( $�L +  ,VR_NO_BUS       1    , -̜ $�L -�  $�L -�  $�\ -̜ $�\ -̜ $�L +  ,VR_NO_BUS       1    , .�( $�L /�h $�L /�h $�\ .�( $�\ .�( $�L +  ,VR_NO_BUS       1    , o0 $�L Q� $�L Q� $�\ o0 $�\ o0 $�L +  ,VR_NO_BUS       1    , �� &�� @ &�� @ &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , �h &�� �� &�� �� &�� �h &�� �h &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , C� &�� _  &�� _  &�� C� &�� C� &�� +  ,VR_NO_BUS       1    , /� &�� 9� &�� 9� &�� /� &�� /� &�� +  ,VR_NO_BUS       1    , �h &�� �� &�� �� &�� �h &�� �h &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , �� &�� �� &�� �� &�� �� &�� �� &�� +  ,VR_NO_BUS       1    , `< $�L j  $�L j  $�\ `< $�\ `< $�L +  ,VR_NO_BUS       1    , ` $�L d  $�L d  $�\ ` $�\ ` $�L +  ,VR_NO_BUS       1    , 4� $�L >� $�L >� $�\ 4� $�\ 4� $�L +  ,VR_NO_BUS       1    , 4� $�L 8� $�L 8� $�\ 4� $�\ 4� $�L +  ,VR_NO_BUS       1    , .� $�L 2� $�L 2� $�\ .� $�\ .� $�L +  ,VR_NO_BUS       1    , (� $�L ,� $�L ,� $�\ (� $�\ (� $�L +  ,VR_NO_BUS       1    , �� $�L � $�L � $�\ �� $�\ �� $�L +  ,VR_NO_BUS       1    , �� $�L � $�L � $�\ �� $�\ �� $�L +  ,VR_NO_BUS       1    , �| $�L �@ $�L �@ $�\ �| $�\ �| $�L +  ,VR_NO_BUS       1    ,  �< $�L  �  $�L  �  $�\  �< $�\  �< $�L +  ,VR_NO_BUS       1    , !� $�L !�  $�L !�  $�\ !� $�\ !� $�L +  ,VR_NO_BUS       1    , "� $�L "�  $�L "�  $�\ "� $�\ "� $�L +  ,VR_NO_BUS       1    , #� $�L #�  $�L #�  $�\ #� $�\ #� $�L +  ,VR_NO_BUS       1    , $u� $�L $� $�L $� $�\ $u� $�\ $u� $�L +  ,VR_NO_BUS       1    , %u� $�L %y� $�L %y� $�\ %u� $�\ %u� $�L +  ,VR_NO_BUS       1    , �X $�L �@ $�L �@ $�\ �X $�\ �X $�L +  ,VR_NO_BUS       1    , �X $�L �@ $�L �@ $�\ �X $�\ �X $�L +  ,VR_NO_BUS       1    , �< $�L �  $�L �  $�\ �< $�\ �< $�L +  ,VR_NO_BUS       1    , � $�L �  $�L �  $�\ � $�\ � $�L +  ,VR_NO_BUS       1    , � $�L #  $�L #  $�\ � $�\ � $�L +  ,VR_NO_BUS       1    ,  $�L   $�L   $�\  $�\  $�L +  ,VR_NO_BUS       1    , �� $�L �� $�L �� $�\ �� $�\ �� $�L +  ,VR_NO_BUS       1    , �� $�L �� $�L �� $�\ �� $�\ �� $�L +  ,VR_NO_BUS       1    , Sh $�L n� $�L n� $�\ Sh $�\ Sh $�L +  ,VR_NO_BUS       1    , d� $�L h� $�L h� $�\ d� $�\ d� $�L +  ,VR_NO_BUS       1    , 9� $�L C� $�L C� $�\ 9� $�\ 9� $�L +  ,VR_NO_BUS       1    , | $�L @ $�L @ $�\ | $�\ | $�L +  ,VR_NO_BUS       1    , X $�L @ $�L @ $�\ X $�\ X $�L +  ,VR_NO_BUS       1    , y� $�L �@ $�L �@ $�\ y� $�\ y� $�L +  ,VR_NO_BUS       1    , s� $�L �@ $�L �@ $�\ s� $�\ s� $�L +  ,VR_NO_BUS       1    , *� "�� *�  "�� *�  "�� *� "�� *� "�� +  ,VR_NO_BUS       1    , +�� "�� +�� "�� +�� "�� +�� "�� +�� "�� +  ,VR_NO_BUS       1    , ,�� "�� ,�� "�� ,�� "�� ,�� "�� ,�� "�� +  ,VR_NO_BUS       1    , -�� "�� /�h "�� /�h "�� -�� "�� -�� "�� +  ,VR_NO_BUS       1    , o0 "�� Q� "�� Q� "�� o0 "�� o0 "�� +  ,VR_NO_BUS       1    , Ҩ $�L �  $�L �  $�\ Ҩ $�\ Ҩ $�L +  ,VR_NO_BUS       1    , � $�L �  $�L �  $�\ � $�\ � $�L +  ,VR_NO_BUS       1    , I� $�L e  $�L e  $�\ I� $�\ I� $�L +  ,VR_NO_BUS       1    , 5� $�L ?� $�L ?� $�\ 5� $�\ 5� $�L +  ,VR_NO_BUS       1    , 5� $�L 9� $�L 9� $�\ 5� $�\ 5� $�L +  ,VR_NO_BUS       1    , /� $�L 3� $�L 3� $�\ /� $�\ /� $�L +  ,VR_NO_BUS       1    , � $�L � $�L � $�\ � $�\ � $�L +  ,VR_NO_BUS       1    , �| $�L �@ $�L �@ $�\ �| $�\ �| $�L +  ,VR_NO_BUS       1    , 	�X $�L 	�@ $�L 	�@ $�\ 	�X $�\ 	�X $�L +  ,VR_NO_BUS       1    , 
�X $�L 
�@ $�L 
�@ $�\ 
�X $�\ 
�X $�L +  ,VR_NO_BUS       1    , � "�� � "�� � "�� � "�� � "�� +  ,VR_NO_BUS       1    , �� "�� � "�� � "�� �� "�� �� "�� +  ,VR_NO_BUS       1    , �| "�� �@ "�� �@ "�� �| "�� �| "�� +  ,VR_NO_BUS       1    ,  �X "��  �@ "��  �@ "��  �X "��  �X "�� +  ,VR_NO_BUS       1    , !�< "�� !�  "�� !�  "�� !�< "�� !�< "�� +  ,VR_NO_BUS       1    , "� "�� "�  "�� "�  "�� "� "�� "� "�� +  ,VR_NO_BUS       1    , #{� "�� #�� "�� #�� "�� #{� "�� #{� "�� +  ,VR_NO_BUS       1    , $V� "�� $`� "�� $`� "�� $V� "�� $V� "�� +  ,VR_NO_BUS       1    , %V� "�� %Z� "�� %Z� "�� %V� "�� %V� "�� +  ,VR_NO_BUS       1    , &+| "�� &5@ "�� &5@ "�� &+| "�� &+| "�� +  ,VR_NO_BUS       1    , &�� "�� &�@ "�� &�@ "�� &�� "�� &�� "�� +  ,VR_NO_BUS       1    , '�X "�� '�@ "�� '�@ "�� '�X "�� '�X "�� +  ,VR_NO_BUS       1    , (�X "�� (�@ "�� (�@ "�� (�X "�� (�X "�� +  ,VR_NO_BUS       1    , )w< "�� )�  "�� )�  "�� )w< "�� )w< "�� +  ,VR_NO_BUS       1    , )� "�� )�  "�� )�  "�� )� "�� )� "�� +  ,VR_NO_BUS       1    , �h "�� �� "�� �� "�� �h "�� �h "�� +  ,VR_NO_BUS       1    , Sh "�� n� "�� n� "�� Sh "�� Sh "�� +  ,VR_NO_BUS       1    , ?� "�� I� "�� I� "�� ?� "�� ?� "�� +  ,VR_NO_BUS       1    , | "�� $@ "�� $@ "�� | "�� | "�� +  ,VR_NO_BUS       1    , X "�� @ "�� @ "�� X "�� X "�� +  ,VR_NO_BUS       1    , X "�� @ "�� @ "�� X "�� X "�� +  ,VR_NO_BUS       1    , y� "�� �@ "�� �@ "�� y� "�� y� "�� +  ,VR_NO_BUS       1    , f< "�� p  "�� p  "�� f< "�� f< "�� +  ,VR_NO_BUS       1    , Ѩ "�� �  "�� �  "�� Ѩ "�� Ѩ "�� +  ,VR_NO_BUS       1    , � "�� �  "�� �  "�� � "�� � "�� +  ,VR_NO_BUS       1    , � "�� �  "�� �  "�� � "�� � "�� +  ,VR_NO_BUS       1    , �� "�� �� "�� �� "�� �� "�� �� "�� +  ,VR_NO_BUS       1    , h "�� 8� "�� 8� "�� h "�� h "�� +  ,VR_NO_BUS       1    , .� "�� 2� "�� 2� "�� .� "�� .� "�� +  ,VR_NO_BUS       1    , � "�� � "�� � "�� � "�� � "�� +  ,VR_NO_BUS       1    , �� "�� �� "�� �� "�� �� "�� �� "�� +  ,VR_NO_BUS       1    , �� "�� �� "�� �� "�� �� "�� �� "�� +  ,VR_NO_BUS       1    , h "�� 3� "�� 3� "�� h "�� h "�� +  ,VR_NO_BUS       1    , )� "�� -� "�� -� "�� )� "�� )� "�� +  ,VR_NO_BUS       1    , 	#� "�� 	'� "�� 	'� "�� 	#� "�� 	#� "�� +  ,VR_NO_BUS       1    , 	�� "�� 
� "�� 
� "�� 	�� "�� 	�� "�� +  ,VR_NO_BUS       1    , 
�� "�� 
�� "�� 
�� "�� 
�� "�� 
�� "�� +  ,VR_NO_BUS       1    , � "�� �� "�� �� "�� � "�� � "�� +  ,VR_NO_BUS       1    , wh "�� �� "�� �� "�� wh "�� wh "�� +  ,VR_NO_BUS       1    , c� "�� m� "�� m� "�� c� "�� c� "�� +  ,VR_NO_BUS       1    , �( "�� � "�� � "�� �( "�� �( "�� +  ,VR_NO_BUS       1    , �� "�� � "�� � "�� �� "�� �� "�� +  ,VR_NO_BUS       1    , ژ "�� ހ "�� ހ "�� ژ "�� ژ "�� +  ,VR_NO_BUS       1    , _h "�� z� "�� z� "�� _h "�� _h "�� +  ,VR_NO_BUS       1    , � "�� 6@ "�� 6@ "�� � "�� � "�� +  ,VR_NO_BUS       1    , %��  � %��  � %��  �$ %��  �$ %��  � +  ,VR_NO_BUS       1    , &Ǽ  � &р  � &р  �$ &Ǽ  �$ &Ǽ  � +  ,VR_NO_BUS       1    , 'ǘ  � 'ˀ  � 'ˀ  �$ 'ǘ  �$ 'ǘ  � +  ,VR_NO_BUS       1    , (�|  � (�@  � (�@  �$ (�|  �$ (�|  � +  ,VR_NO_BUS       1    , )�X  � )�@  � )�@  �$ )�X  �$ )�X  � +  ,VR_NO_BUS       1    , *q<  � *{   � *{   �$ *q<  �$ *q<  � +  ,VR_NO_BUS       1    , +q  � +u   � +u   �$ +q  �$ +q  � +  ,VR_NO_BUS       1    , ,k  � ,o   � ,o   �$ ,k  �$ ,k  � +  ,VR_NO_BUS       1    , -?�  � -I�  � -I�  �$ -?�  �$ -?�  � +  ,VR_NO_BUS       1    , .�  � .$�  � .$�  �$ .�  �$ .�  � +  ,VR_NO_BUS       1    , .�(  � /�h  � /�h  �$ .�(  �$ .�(  � +  ,VR_NO_BUS       1    , o0  � Q�  � Q�  �$ o0  �$ o0  � +  ,VR_NO_BUS       1    , G� "�� K� "�� K� "�� G� "�� G� "�� +  ,VR_NO_BUS       1    , �� "�� @ "�� @ "�� �� "�� �� "�� +  ,VR_NO_BUS       1    , �h "�� �� "�� �� "�� �h "�� �h "�� +  ,VR_NO_BUS       1    , @�  � J�  � J�  �$ @�  �$ @�  � +  ,VR_NO_BUS       1    , @�  � D�  � D�  �$ @�  �$ @�  � +  ,VR_NO_BUS       1    , :�  � >�  � >�  �$ :�  �$ :�  � +  ,VR_NO_BUS       1    , �  � �  � �  �$ �  �$ �  � +  ,VR_NO_BUS       1    , �  � �  � �  �$ �  �$ �  � +  ,VR_NO_BUS       1    , 	�  � �  � �  �$ 	�  �$ 	�  � +  ,VR_NO_BUS       1    , o(  � ��  � ��  �$ o(  �$ o(  � +  ,VR_NO_BUS       1    , [|  � e@  � e@  �$ [|  �$ [|  � +  ,VR_NO_BUS       1    , [X  � _@  � _@  �$ [X  �$ [X  � +  ,VR_NO_BUS       1    ,  0<  �  :   �  :   �$  0<  �$  0<  � +  ,VR_NO_BUS       1    , !0  � !4   � !4   �$ !0  �$ !0  � +  ,VR_NO_BUS       1    , "*  � ".   � ".   �$ "*  �$ "*  � +  ,VR_NO_BUS       1    , #$  � #(   � #(   �$ #$  �$ #$  � +  ,VR_NO_BUS       1    , #��  � $�  � $�  �$ #��  �$ #��  � +  ,VR_NO_BUS       1    , $��  � $��  � $��  �$ $��  �$ $��  � +  ,VR_NO_BUS       1    , u�  � y�  � y�  �$ u�  �$ u�  � +  ,VR_NO_BUS       1    , �  � 5   � 5   �$ �  �$ �  � +  ,VR_NO_BUS       1    , +  � /   � /   �$ +  �$ +  � +  ,VR_NO_BUS       1    , �(  � �  � �  �$ �(  �$ �(  � +  ,VR_NO_BUS       1    , ��  � �  � �  �$ ��  �$ ��  � +  ,VR_NO_BUS       1    , �|  � �@  � �@  �$ �|  �$ �|  � +  ,VR_NO_BUS       1    , �X  � �@  � �@  �$ �X  �$ �X  � +  ,VR_NO_BUS       1    , �<  � �   � �   �$ �<  �$ �<  � +  ,VR_NO_BUS       1    , �  � �   � �   �$ �  �$ �  � +  ,VR_NO_BUS       1    , �  � *@  � *@  �$ �  �$ �  � +  ,VR_NO_BUS       1    , ��  � �@  � �@  �$ ��  �$ ��  � +  ,VR_NO_BUS       1    , �X  � �@  � �@  �$ �X  �$ �X  � +  ,VR_NO_BUS       1    , r<  � |   � |   �$ r<  �$ r<  � +  ,VR_NO_BUS       1    , r  � v   � v   �$ r  �$ r  � +  ,VR_NO_BUS       1    , l  � p   � p   �$ l  �$ l  � +  ,VR_NO_BUS       1    , *�  � *�   � *�  G� *� G� *�  � +  ,VR_NO_BUS       1    , +��  � +��  � +�� G� +�� G� +��  � +  ,VR_NO_BUS       1    , ,��  � ,��  � ,�� G� ,�� G� ,��  � +  ,VR_NO_BUS       1    , -��  � -��  � -�� G� -�� G� -��  � +  ,VR_NO_BUS       1    , .��  � /�h  � /�h G� .�� G� .��  � +  ,VR_NO_BUS       1    , o0  � Q�  � Q� G� o0 G� o0  � +  ,VR_NO_BUS       1    , G�  � K�  � K�  �$ G�  �$ G�  � +  ,VR_NO_BUS       1    , �h  � ��  � ��  �$ �h  �$ �h  � +  ,VR_NO_BUS       1    , ��  � ��  � ��  �$ ��  �$ ��  � +  ,VR_NO_BUS       1    , ��  � ��  � ��  �$ ��  �$ ��  � +  ,VR_NO_BUS       1    , ��  � ��  � ��  �$ ��  �$ ��  � +  ,VR_NO_BUS       1    , ��  � ��  � ��  �$ ��  �$ ��  � +  ,VR_NO_BUS       1    , ��  � ��  � ��  �$ ��  �$ ��  � +  ,VR_NO_BUS       1    , 	��  � 	��  � 	��  �$ 	��  �$ 	��  � +  ,VR_NO_BUS       1    , 
{�  � 
�  � 
�  �$ 
{�  �$ 
{�  � +  ,VR_NO_BUS       1    , a|  � k@  � k@ G� a| G� a|  � +  ,VR_NO_BUS       1    , aX  � e@  � e@ G� aX G� aX  � +  ,VR_NO_BUS       1    , [X  � _@  � _@ G� [X G� [X  � +  ,VR_NO_BUS       1    , ��  � �@  � �@ G� �� G� ��  � +  ,VR_NO_BUS       1    ,  �X  �  �@  �  �@ G�  �X G�  �X  � +  ,VR_NO_BUS       1    , !�<  � !�   � !�  G� !�< G� !�<  � +  ,VR_NO_BUS       1    , "��  � "��  � "�� G� "�� G� "��  � +  ,VR_NO_BUS       1    , #��  � #��  � #�� G� #�� G� #��  � +  ,VR_NO_BUS       1    , ${�  � $�  � $� G� ${� G� ${�  � +  ,VR_NO_BUS       1    , %P�  � %Z�  � %Z� G� %P� G� %P�  � +  ,VR_NO_BUS       1    , &P�  � &T�  � &T� G� &P� G� &P�  � +  ,VR_NO_BUS       1    , '%|  � '/@  � '/@ G� '%| G� '%|  � +  ,VR_NO_BUS       1    , (%X  � ()@  � ()@ G� (%X G� (%X  � +  ,VR_NO_BUS       1    , )X  � )#@  � )#@ G� )X G� )X  � +  ,VR_NO_BUS       1    , )�<  � )�   � )�  G� )�< G� )�<  � +  ,VR_NO_BUS       1    , �X  � �@  � �@ G� �X G� �X  � +  ,VR_NO_BUS       1    , �  � 6@  � 6@ G� � G� �  � +  ,VR_NO_BUS       1    , ,X  � 0@  � 0@ G� ,X G� ,X  � +  ,VR_NO_BUS       1    , &X  � *@  � *@ G� &X G� &X  � +  ,VR_NO_BUS       1    ,  X  � $@  � $@ G�  X G�  X  � +  ,VR_NO_BUS       1    , �<  � �   � �  G� �< G� �<  � +  ,VR_NO_BUS       1    , �  � �   � �  G� � G� �  � +  ,VR_NO_BUS       1    , ��  � ��  � �� G� �� G� ��  � +  ,VR_NO_BUS       1    , 5h  � P�  � P� G� 5h G� 5h  � +  ,VR_NO_BUS       1    , F�  � J�  � J� G� F� G� F�  � +  ,VR_NO_BUS       1    , @�  � D�  � D� G� @� G� @�  � +  ,VR_NO_BUS       1    , �  � �  � � G� � G� �  � +  ,VR_NO_BUS       1    , �(  � ��  � �� G� �( G� �(  � +  ,VR_NO_BUS       1    , ��  � ��  � �� G� �� G� ��  � +  ,VR_NO_BUS       1    , ��  � ��  � �� G� �� G� ��  � +  ,VR_NO_BUS       1    , ��  � ��  � �� G� �� G� ��  � +  ,VR_NO_BUS       1    , ��  � ��  � �� G� �� G� ��  � +  ,VR_NO_BUS       1    , C�  � _   � _  G� C� G� C�  � +  ,VR_NO_BUS       1    , U  � Y   � Y  G� U G� U  � +  ,VR_NO_BUS       1    , �(  � �  � � G� �( G� �(  � +  ,VR_NO_BUS       1    , ��  � �   � �  G� �� G� ��  � +  ,VR_NO_BUS       1    , �  � �   � �  G� � G� �  � +  ,VR_NO_BUS       1    , 	��  � 	��  � 	�� G� 	�� G� 	��  � +  ,VR_NO_BUS       1    , 
��  � 
��  � 
�� G� 
�� G� 
��  � +  ,VR_NO_BUS       1    , o�  � y�  � y� G� o� G� o�  � +  ,VR_NO_BUS       1    , o�  � s�  � s� G� o� G� o�  � +  ,VR_NO_BUS       1    , �(  � ��  � �� G� �( G� �(  � +  ,VR_NO_BUS       1    , �  � �  � � G� � G� �  � +  ,VR_NO_BUS       1    , ��  � �  � � G� �� G� ��  � +  ,VR_NO_BUS       1    , �|  � �@  � �@ G� �| G� �|  � +  ,VR_NO_BUS       1    , $E( � $`� � $`� � $E( � $E( � +  ,VR_NO_BUS       1    , %1| � %;@ � %;@ � %1| � %1| � +  ,VR_NO_BUS       1    , &1X � &5@ � &5@ � &1X � &1X � +  ,VR_NO_BUS       1    , '+X � '/@ � '/@ � '+X � '+X � +  ,VR_NO_BUS       1    , '� � (
  � (
  � '� � '� � +  ,VR_NO_BUS       1    , (k� � (�  � (�  � (k� � (k� � +  ,VR_NO_BUS       1    , )} � )�  � )�  � )} � )} � +  ,VR_NO_BUS       1    , *w � *{  � *{  � *w � *w � +  ,VR_NO_BUS       1    , +K� � +U� � +U� � +K� � +K� � +  ,VR_NO_BUS       1    , ,K� � ,O� � ,O� � ,K� � ,K� � +  ,VR_NO_BUS       1    , - � � -*� � -*� � - � � - � � +  ,VR_NO_BUS       1    , -�( � -�� � -�� � -�( � -�( � +  ,VR_NO_BUS       1    , .�� � /�h � /�h � .�� � .�� � +  ,VR_NO_BUS       1    , o0 � Q� � Q� � o0 � o0 � +  ,VR_NO_BUS       1    , �h  � ��  � �� G� �h G� �h  � +  ,VR_NO_BUS       1    , L� � P� � P� � L� � L� � +  ,VR_NO_BUS       1    , !� � +� � +� � !� � !� � +  ,VR_NO_BUS       1    , !� � %� � %� � !� � !� � +  ,VR_NO_BUS       1    , � � � � � � � � � � +  ,VR_NO_BUS       1    , �| � �@ � �@ � �| � �| � +  ,VR_NO_BUS       1    , [� � w@ � w@ � [� � [� � +  ,VR_NO_BUS       1    , H< � R  � R  � H< � H< � +  ,VR_NO_BUS       1    , H � L  � L  � H � H � +  ,VR_NO_BUS       1    , B � F  � F  � B � B � +  ,VR_NO_BUS       1    , � �  � �  � � � � � � +  ,VR_NO_BUS       1    , � � �� � �� � � � � � +  ,VR_NO_BUS       1    ,  � �  �� �  �� �  � �  � � +  ,VR_NO_BUS       1    , !� � !� � !� � !� � !� � +  ,VR_NO_BUS       1    , "� � "� � "� � "� � "� � +  ,VR_NO_BUS       1    , #ߘ � #� � #� � #ߘ � #ߘ � +  ,VR_NO_BUS       1    , 
�� � 
�� � 
�� � 
�� � 
�� � +  ,VR_NO_BUS       1    , ^( � y� � y� � ^( � ^( � +  ,VR_NO_BUS       1    , J| � T@ � T@ � J| � J| � +  ,VR_NO_BUS       1    , %< � /  � /  � %< � %< � +  ,VR_NO_BUS       1    , % � )  � )  � % � % � +  ,VR_NO_BUS       1    , �� � � � � � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �@ � �@ � �� � �� � +  ,VR_NO_BUS       1    , �X � �@ � �@ � �X � �X � +  ,VR_NO_BUS       1    , �< � �  � �  � �< � �< � +  ,VR_NO_BUS       1    , � �   �   � � � � � +  ,VR_NO_BUS       1    ,  �   �   �  �  � +  ,VR_NO_BUS       1    , f� � �  � �  � f� � f� � +  ,VR_NO_BUS       1    , R� � \� � \� � R� � R� � +  ,VR_NO_BUS       1    , R� � V� � V� � R� � R� � +  ,VR_NO_BUS       1    , *�X �� *�@ �� *�@ �� *�X �� *�X �� +  ,VR_NO_BUS       1    , +�X �� +�@ �� +�@ �� +�X �� +�X �� +  ,VR_NO_BUS       1    , ,S� �� ,o  �� ,o  �� ,S� �� ,S� �� +  ,VR_NO_BUS       1    , -e �� -i  �� -i  �� -e �� -e �� +  ,VR_NO_BUS       1    , -ʨ �� /�h �� /�h �� -ʨ �� -ʨ �� +  ,VR_NO_BUS       1    , o0 �� Q� �� Q� �� o0 �� o0 �� +  ,VR_NO_BUS       1    , "� � ,� � ,� � "� � "� � +  ,VR_NO_BUS       1    , "� � &� � &� � "� � "� � +  ,VR_NO_BUS       1    , � �  � �  � � � � � � +  ,VR_NO_BUS       1    , �� � �  � �  � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , 	h � 	'� � 	'� � 	h � 	h � +  ,VR_NO_BUS       1    , 	�� � 
� � 
� � 	�� � 	�� � +  ,VR_NO_BUS       1    , gX �� k@ �� k@ �� gX �� gX �� +  ,VR_NO_BUS       1    , aX �� e@ �� e@ �� aX �� aX �� +  ,VR_NO_BUS       1    , [X �� _@ �� _@ �� [X �� [X �� +  ,VR_NO_BUS       1    , �� �� �@ �� �@ �� �� �� �� �� +  ,VR_NO_BUS       1    ,  �X ��  �@ ��  �@ ��  �X ��  �X �� +  ,VR_NO_BUS       1    , !�< �� !�  �� !�  �� !�< �� !�< �� +  ,VR_NO_BUS       1    , "� �� "�  �� "�  �� "� �� "� �� +  ,VR_NO_BUS       1    , #{� �� #�� �� #�� �� #{� �� #{� �� +  ,VR_NO_BUS       1    , ${� �� $� �� $� �� ${� �� ${� �� +  ,VR_NO_BUS       1    , %u� �� %y� �� %y� �� %u� �� %u� �� +  ,VR_NO_BUS       1    , %�h �� %�� �� %�� �� %�h �� %�h �� +  ,VR_NO_BUS       1    , &Ǽ �� &р �� &р �� &Ǽ �� &Ǽ �� +  ,VR_NO_BUS       1    , 'ǘ �� 'ˀ �� 'ˀ �� 'ǘ �� 'ǘ �� +  ,VR_NO_BUS       1    , (�� �� (ŀ �� (ŀ �� (�� �� (�� �� +  ,VR_NO_BUS       1    , )�| �� )�@ �� )�@ �� )�| �� )�| �� +  ,VR_NO_BUS       1    , ]� �� a� �� a� �� ]� �� ]� �� +  ,VR_NO_BUS       1    , 2| �� <@ �� <@ �� 2| �� 2| �� +  ,VR_NO_BUS       1    , 2X �� 6@ �� 6@ �� 2X �� 2X �� +  ,VR_NO_BUS       1    , ,X �� 0@ �� 0@ �� ,X �� ,X �� +  ,VR_NO_BUS       1    , < ��   ��   �� < �� < �� +  ,VR_NO_BUS       1    ,  ��   ��   ��  ��  �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , g| �� q@ �� q@ �� g| �� g| �� +  ,VR_NO_BUS       1    , o0 � Q� � Q� � o0 � o0 � +  ,VR_NO_BUS       1    , G� �� K� �� K� �� G� �� G� �� +  ,VR_NO_BUS       1    , �� �� @ �� @ �� �� �� �� �� +  ,VR_NO_BUS       1    , �X �� @ �� @ �� �X �� �X �� +  ,VR_NO_BUS       1    , �X �� �@ �� �@ �� �X �� �X �� +  ,VR_NO_BUS       1    , �< �� �  �� �  �� �< �� �< �� +  ,VR_NO_BUS       1    , 7� �� S  �� S  �� 7� �� 7� �� +  ,VR_NO_BUS       1    , I �� M  �� M  �� I �� I �� +  ,VR_NO_BUS       1    , �� �� �  �� �  �� �� �� �� �� +  ,VR_NO_BUS       1    , 	�� �� 	�� �� 	�� �� 	�� �� 	�� �� +  ,VR_NO_BUS       1    , 
�� �� 
�� �� 
�� �� 
�� �� 
�� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , �� �� �� �� �� �� �� �� �� �� +  ,VR_NO_BUS       1    , ]� �� g� �� g� �� ]� �� ]� �� +  ,VR_NO_BUS       1    , !� � !�  � !�  � !� � !� � +  ,VR_NO_BUS       1    , "�� � "�� � "�� � "�� � "�� � +  ,VR_NO_BUS       1    , #�� � #�� � #�� � #�� � #�� � +  ,VR_NO_BUS       1    , ${� � $� � $� � ${� � ${� � +  ,VR_NO_BUS       1    , %P� � %Z� � %Z� � %P� � %P� � +  ,VR_NO_BUS       1    , &P� � &T� � &T� � &P� � &P� � +  ,VR_NO_BUS       1    , 'J� � 'N� � 'N� � 'J� � 'J� � +  ,VR_NO_BUS       1    , (| � ()@ � ()@ � (| � (| � +  ,VR_NO_BUS       1    , )X � )#@ � )#@ � )X � )X � +  ,VR_NO_BUS       1    , *X � *@ � *@ � *X � *X � +  ,VR_NO_BUS       1    , *�< � *�  � *�  � *�< � *�< � +  ,VR_NO_BUS       1    , +� � ,O� � ,O� � +� � +� � +  ,VR_NO_BUS       1    , ,�h � ,�� � ,�� � ,�h � ,�h � +  ,VR_NO_BUS       1    , -�h � -�� � -�� � -�h � -�h � +  ,VR_NO_BUS       1    , .�� � /�h � /�h � .�� � .�� � +  ,VR_NO_BUS       1    , (( � C� � C� � (( � (( � +  ,VR_NO_BUS       1    , | � @ � @ � | � | � +  ,VR_NO_BUS       1    , X � @ � @ � X � X � +  ,VR_NO_BUS       1    , X � @ � @ � X � X � +  ,VR_NO_BUS       1    , X � @ � @ � X � X � +  ,VR_NO_BUS       1    , �< � �  � �  � �< � �< � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �( � � � � � �( � �( � +  ,VR_NO_BUS       1    , �| � �@ � �@ � �| � �| � +  ,VR_NO_BUS       1    , �X � �@ � �@ � �X � �X � +  ,VR_NO_BUS       1    , �X � �@ � �@ � �X � �X � +  ,VR_NO_BUS       1    , �< � �  � �  � �< � �< � +  ,VR_NO_BUS       1    ,  � �  �  �  �  �  � �  � � +  ,VR_NO_BUS       1    , 	#� � 	'� � 	'� � 	#� � 	#� � +  ,VR_NO_BUS       1    , 	�� � 	�  � 	�  � 	�� � 	�� � +  ,VR_NO_BUS       1    , 
d( � 
� � 
� � 
d( � 
d( � +  ,VR_NO_BUS       1    , P| � Z@ � Z@ � P| � P| � +  ,VR_NO_BUS       1    , �� � �@ � �@ � �� � �� � +  ,VR_NO_BUS       1    , 8� � T@ � T@ � 8� � 8� � +  ,VR_NO_BUS       1    , %< � /  � /  � %< � %< � +  ,VR_NO_BUS       1    , �� � �  � �  � �� � �� � +  ,VR_NO_BUS       1    , � � �  � �  � � � � � +  ,VR_NO_BUS       1    , � � �  � �  � � � � � +  ,VR_NO_BUS       1    , � � �  � �  � � � � � +  ,VR_NO_BUS       1    , j� � t� � t� � j� � j� � +  ,VR_NO_BUS       1    , �h � �� � �� � �h � �h � +  ,VR_NO_BUS       1    , ¼ � ̀ � ̀ � ¼ � ¼ � +  ,VR_NO_BUS       1    ,  � ƀ � ƀ �  �  � +  ,VR_NO_BUS       1    , *@h r< *[� r< *[� �L *@h �L *@h r< +  ,VR_NO_BUS       1    , +Q� r< +U� r< +U� �L +Q� �L +Q� r< +  ,VR_NO_BUS       1    , ,&� r< ,0� r< ,0� �L ,&� �L ,&� r< +  ,VR_NO_BUS       1    , -&� r< -*� r< -*� �L -&� �L -&� r< +  ,VR_NO_BUS       1    , -ʨ r< -�  r< -�  �L -ʨ �L -ʨ r< +  ,VR_NO_BUS       1    , .f� r< /�h r< /�h �L .f� �L .f� r< +  ,VR_NO_BUS       1    , o0 r< Q� r< Q� �L o0 �L o0 r< +  ,VR_NO_BUS       1    , Ҩ � �  � �  � Ҩ � Ҩ � +  ,VR_NO_BUS       1    , �( � �� � �� � �( � �( � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , ( �  � �  � � ( � ( � +  ,VR_NO_BUS       1    , �� � �  � �  � �� � �� � +  ,VR_NO_BUS       1    , � � �  � �  � � � � � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , h � -� � -� � h � h � +  ,VR_NO_BUS       1    , �� r< �� r< �� �L �� �L �� r< +  ,VR_NO_BUS       1    , z� r< �� r< �� �L z� �L z� r< +  ,VR_NO_BUS       1    , z� r< ~� r< ~� �L z� �L z� r< +  ,VR_NO_BUS       1    ,  O| r<  Y@ r<  Y@ �L  O| �L  O| r< +  ,VR_NO_BUS       1    ,  �� r<  �@ r<  �@ �L  �� �L  �� r< +  ,VR_NO_BUS       1    , !�X r< !�@ r< !�@ �L !�X �L !�X r< +  ,VR_NO_BUS       1    , "�X r< "�@ r< "�@ �L "�X �L "�X r< +  ,VR_NO_BUS       1    , #�X r< #�@ r< #�@ �L #�X �L #�X r< +  ,VR_NO_BUS       1    , $�� r< $�@ r< $�@ �L $�� �L $�� r< +  ,VR_NO_BUS       1    , %� r< %;@ r< %;@ �L %� �L %� r< +  ,VR_NO_BUS       1    , &1X r< &5@ r< &5@ �L &1X �L &1X r< +  ,VR_NO_BUS       1    , '+X r< '/@ r< '/@ �L '+X �L '+X r< +  ,VR_NO_BUS       1    , ( < r< (
  r< (
  �L ( < �L ( < r< +  ,VR_NO_BUS       1    , (�( r< (ŀ r< (ŀ �L (�( �L (�( r< +  ,VR_NO_BUS       1    , )�� r< )�� r< )�� �L )�� �L )�� r< +  ,VR_NO_BUS       1    ,  r<   r<   �L  �L  r< +  ,VR_NO_BUS       1    , �� r< �� r< �� �L �� �L �� r< +  ,VR_NO_BUS       1    , �� r< �� r< �� �L �� �L �� r< +  ,VR_NO_BUS       1    , Sh r< n� r< n� �L Sh �L Sh r< +  ,VR_NO_BUS       1    , d� r< h� r< h� �L d� �L d� r< +  ,VR_NO_BUS       1    , 9� r< C� r< C� �L 9� �L 9� r< +  ,VR_NO_BUS       1    , 9� r< =� r< =� �L 9� �L 9� r< +  ,VR_NO_BUS       1    , | r< @ r< @ �L | �L | r< +  ,VR_NO_BUS       1    , X r< @ r< @ �L X �L X r< +  ,VR_NO_BUS       1    , �< r< �  r< �  �L �< �L �< r< +  ,VR_NO_BUS       1    , � r< �  r< �  �L � �L � r< +  ,VR_NO_BUS       1    , � r< �  r< �  �L � �L � r< +  ,VR_NO_BUS       1    , � r< �  r< �  �L � �L � r< +  ,VR_NO_BUS       1    , �� r< �� r< �� �L �� �L �� r< +  ,VR_NO_BUS       1    , �� r< �� r< �� �L �� �L �� r< +  ,VR_NO_BUS       1    , �� r< �� r< �� �L �� �L �� r< +  ,VR_NO_BUS       1    , *h r< E� r< E� �L *h �L *h r< +  ,VR_NO_BUS       1    , � r<  � r<  � �L � �L � r< +  ,VR_NO_BUS       1    , � r< � r< � �L � �L � r< +  ,VR_NO_BUS       1    , |( r< �� r< �� �L |( �L |( r< +  ,VR_NO_BUS       1    , �� r< �� r< �� �L �� �L �� r< +  ,VR_NO_BUS       1    , b| r< l@ r< l@ �L b| �L b| r< +  ,VR_NO_BUS       1    , 	bX r< 	f@ r< 	f@ �L 	bX �L 	bX r< +  ,VR_NO_BUS       1    , 
7< r< 
A  r< 
A  �L 
7< �L 
7< r< +  ,VR_NO_BUS       1    , 7 r< ;  r< ;  �L 7 �L 7 r< +  ,VR_NO_BUS       1    , � r< � r< � �L � �L � r< +  ,VR_NO_BUS       1    , � r< �� r< �� �L � �L � r< +  ,VR_NO_BUS       1    , R( r< m� r< m� �L R( �L R( r< +  ,VR_NO_BUS       1    , >| r< H@ r< H@ �L >| �L >| r< +  ,VR_NO_BUS       1    , � r< #  r< #  �L � �L � r< +  ,VR_NO_BUS       1    , $� Kt $"  Kt $"  r� $� r� $� Kt +  ,VR_NO_BUS       1    , % � Kt %  Kt %  r� % � r� % � Kt +  ,VR_NO_BUS       1    , %�� Kt %�@ Kt %�@ r� %�� r� %�� Kt +  ,VR_NO_BUS       1    , &Xh Kt &s� Kt &s� r� &Xh r� &Xh Kt +  ,VR_NO_BUS       1    , 'i� Kt 'm� Kt 'm� r� 'i� r� 'i� Kt +  ,VR_NO_BUS       1    , (>� Kt (H� Kt (H� r� (>� r� (>� Kt +  ,VR_NO_BUS       1    , )>� Kt )B� Kt )B� r� )>� r� )>� Kt +  ,VR_NO_BUS       1    , *| Kt *@ Kt *@ r� *| r� *| Kt +  ,VR_NO_BUS       1    , *�� Kt +@ Kt +@ r� *�� r� *�� Kt +  ,VR_NO_BUS       1    , ,X Kt ,@ Kt ,@ r� ,X r� ,X Kt +  ,VR_NO_BUS       1    , ,�� Kt -@ Kt -@ r� ,�� r� ,�� Kt +  ,VR_NO_BUS       1    , -l� Kt -�@ Kt -�@ r� -l� r� -l� Kt +  ,VR_NO_BUS       1    , .~X Kt /�h Kt /�h r� .~X r� .~X Kt +  ,VR_NO_BUS       1    , o0 Kt Q� Kt Q� r� o0 r� o0 Kt +  ,VR_NO_BUS       1    , �h r< �� r< �� �L �h �L �h r< +  ,VR_NO_BUS       1    , l Kt p  Kt p  r� l r� l Kt +  ,VR_NO_BUS       1    , Ѩ Kt �  Kt �  r� Ѩ r� Ѩ Kt +  ,VR_NO_BUS       1    , � Kt �  Kt �  r� � r� � Kt +  ,VR_NO_BUS       1    , � Kt �  Kt �  r� � r� � Kt +  ,VR_NO_BUS       1    , � Kt �  Kt �  r� � r� � Kt +  ,VR_NO_BUS       1    , �� Kt �� Kt �� r� �� r� �� Kt +  ,VR_NO_BUS       1    , �h Kt �� Kt �� r� �h r� �h Kt +  ,VR_NO_BUS       1    , �� Kt �� Kt �� r� �� r� �� Kt +  ,VR_NO_BUS       1    , z� Kt �� Kt �� r� z� r� z� Kt +  ,VR_NO_BUS       1    , z� Kt ~� Kt ~� r� z� r� z� Kt +  ,VR_NO_BUS       1    ,  t� Kt  x� Kt  x� r�  t� r�  t� Kt +  ,VR_NO_BUS       1    , !n� Kt !r� Kt !r� r� !n� r� !n� Kt +  ,VR_NO_BUS       1    , "C| Kt "M@ Kt "M@ r� "C| r� "C| Kt +  ,VR_NO_BUS       1    , "�� Kt "�@ Kt "�@ r� "�� r� "�� Kt +  ,VR_NO_BUS       1    , #�< Kt #�  Kt #�  r� #�< r� #�< Kt +  ,VR_NO_BUS       1    , 
u� Kt 
� Kt 
� r� 
u� r� 
u� Kt +  ,VR_NO_BUS       1    , u� Kt y� Kt y� r� u� r� u� Kt +  ,VR_NO_BUS       1    , 8� Kt T@ Kt T@ r� 8� r� 8� Kt +  ,VR_NO_BUS       1    , JX Kt N@ Kt N@ r� JX r� JX Kt +  ,VR_NO_BUS       1    , DX Kt H@ Kt H@ r� DX r� DX Kt +  ,VR_NO_BUS       1    , �� Kt �@ Kt �@ r� �� r� �� Kt +  ,VR_NO_BUS       1    , �< Kt �  Kt �  r� �< r� �< Kt +  ,VR_NO_BUS       1    , � Kt �  Kt �  r� � r� � Kt +  ,VR_NO_BUS       1    , �� Kt   Kt   r� �� r� �� Kt +  ,VR_NO_BUS       1    ,  Kt   Kt   r�  r�  Kt +  ,VR_NO_BUS       1    , �� Kt �� Kt �� r� �� r� �� Kt +  ,VR_NO_BUS       1    , �� Kt �@ Kt �@ r� �� r� �� Kt +  ,VR_NO_BUS       1    , �X Kt �@ Kt �@ r� �X r� �X Kt +  ,VR_NO_BUS       1    , r< Kt |  Kt |  r� r< r� r< Kt +  ,VR_NO_BUS       1    , r Kt v  Kt v  r� r r� r Kt +  ,VR_NO_BUS       1    , *~� $� *�@ $� *�@ K� *~� K� *~� $� +  ,VR_NO_BUS       1    , +�X $� +�@ $� +�@ K� +�X K� +�X $� +  ,VR_NO_BUS       1    , +�� $� ,@ $� ,@ K� +�� K� +�� $� +  ,VR_NO_BUS       1    , ,Ш $� ,�  $� ,�  K� ,Ш K� ,Ш $� +  ,VR_NO_BUS       1    , -� $� /�h $� /�h K� -� K� -� $� +  ,VR_NO_BUS       1    , o0 $� Q� $� Q� K� o0 K� o0 $� +  ,VR_NO_BUS       1    , "� Kt ,� Kt ,� r� "� r� "� Kt +  ,VR_NO_BUS       1    , �( Kt �� Kt �� r� �( r� �( Kt +  ,VR_NO_BUS       1    , �� Kt �� Kt �� r� �� r� �� Kt +  ,VR_NO_BUS       1    , t| Kt ~@ Kt ~@ r� t| r� t| Kt +  ,VR_NO_BUS       1    , �� Kt �@ Kt �@ r� �� r� �� Kt +  ,VR_NO_BUS       1    , �< Kt �  Kt �  r� �< r� �< Kt +  ,VR_NO_BUS       1    , �� Kt �� Kt �� r� �� r� �� Kt +  ,VR_NO_BUS       1    , �� Kt �� Kt �� r� �� r� �� Kt +  ,VR_NO_BUS       1    , 	�� Kt 	�� Kt 	�� r� 	�� r� 	�� Kt +  ,VR_NO_BUS       1    , $� $� @  $� @  K� $� K� $� $� +  ,VR_NO_BUS       1    ,  � $�  � $�  � K�  � K�  � $� +  ,VR_NO_BUS       1    ,  |h $�  �� $�  �� K�  |h K�  |h $� +  ,VR_NO_BUS       1    , !�� $� !�� $� !�� K� !�� K� !�� $� +  ,VR_NO_BUS       1    , "b� $� "l� $� "l� K� "b� K� "b� $� +  ,VR_NO_BUS       1    , "�( $� "� $� "� K� "�( K� "�( $� +  ,VR_NO_BUS       1    , #ߘ $� #� $� #� K� #ߘ K� #ߘ $� +  ,VR_NO_BUS       1    , $٘ $� $݀ $� $݀ K� $٘ K� $٘ $� +  ,VR_NO_BUS       1    , %?( $� %Z� $� %Z� K� %?( K� %?( $� +  ,VR_NO_BUS       1    , &9( $� &T� $� &T� K� &9( K� &9( $� +  ,VR_NO_BUS       1    , 'J� $� 'N� $� 'N� K� 'J� K� 'J� $� +  ,VR_NO_BUS       1    , '� $� (
  $� (
  K� '� K� '� $� +  ,VR_NO_BUS       1    , (�( $� (ŀ $� (ŀ K� (�( K� (�( $� +  ,VR_NO_BUS       1    , )e� $� )�  $� )�  K� )e� K� )e� $� +  ,VR_NO_BUS       1    , *� $� *@ $� *@ K� *� K� *� $� +  ,VR_NO_BUS       1    ,  $�   $�   K�  K�  $� +  ,VR_NO_BUS       1    , �� $� �� $� �� K� �� K� �� $� +  ,VR_NO_BUS       1    , �� $� �@ $� �@ K� �� K� �� $� +  ,VR_NO_BUS       1    , x< $� �  $� �  K� x< K� x< $� +  ,VR_NO_BUS       1    , x $� |  $� |  K� x K� x $� +  ,VR_NO_BUS       1    , L� $� V� $� V� K� L� K� L� $� +  ,VR_NO_BUS       1    , L� $� P� $� P� K� L� K� L� $� +  ,VR_NO_BUS       1    , !� $� +� $� +� K� !� K� !� $� +  ,VR_NO_BUS       1    , !� $� %� $� %� K� !� K� !� $� +  ,VR_NO_BUS       1    , �| $�  @ $�  @ K� �| K� �| $� +  ,VR_NO_BUS       1    , �X $� �@ $� �@ K� �X K� �X $� +  ,VR_NO_BUS       1    , �X $� �@ $� �@ K� �X K� �X $� +  ,VR_NO_BUS       1    , U� $� q@ $� q@ K� U� K� U� $� +  ,VR_NO_BUS       1    , gX $� k@ $� k@ K� gX K� gX $� +  ,VR_NO_BUS       1    , aX $� e@ $� e@ K� aX K� aX $� +  ,VR_NO_BUS       1    , "� $� &� $� &� K� "� K� "� $� +  ,VR_NO_BUS       1    , �| $� @ $� @ K� �| K� �| $� +  ,VR_NO_BUS       1    , �X $� �@ $� �@ K� �X K� �X $� +  ,VR_NO_BUS       1    , �< $� �  $� �  K� �< K� �< $� +  ,VR_NO_BUS       1    , � $� �  $� �  K� � K� � $� +  ,VR_NO_BUS       1    , �� $� �� $� �� K� �� K� �� $� +  ,VR_NO_BUS       1    , 	�� $� 	�� $� 	�� K� 	�� K� 	�� $� +  ,VR_NO_BUS       1    , 
�� $� 
�� $� 
�� K� 
�� K� 
�� $� +  ,VR_NO_BUS       1    , o� $� y� $� y� K� o� K� o� $� +  ,VR_NO_BUS       1    , o� $� s� $� s� K� o� K� o� $� +  ,VR_NO_BUS       1    , i� $� m� $� m� K� i� K� i� $� +  ,VR_NO_BUS       1    , >| $� H@ $� H@ K� >| K� >| $� +  ,VR_NO_BUS       1    , >X $� B@ $� B@ K� >X K� >X $� +  ,VR_NO_BUS       1    , < $�   $�   K� < K� < $� +  ,VR_NO_BUS       1    ,  $�   $�   K�  K�  $� +  ,VR_NO_BUS       1    , #�h ܰ $� ܰ $� � #�h � #�h ܰ +  ,VR_NO_BUS       1    , $�� ܰ $�  ܰ $�  � $�� � $�� ܰ +  ,VR_NO_BUS       1    , %� ܰ %�  ܰ %�  � %� � %� ܰ +  ,VR_NO_BUS       1    , &i� ܰ &s� ܰ &s� � &i� � &i� ܰ +  ,VR_NO_BUS       1    , 'i� ܰ 'm� ܰ 'm� � 'i� � 'i� ܰ +  ,VR_NO_BUS       1    , '� ܰ (
  ܰ (
  � '� � '� ܰ +  ,VR_NO_BUS       1    , )  ܰ )  ܰ )  � )  � )  ܰ +  ,VR_NO_BUS       1    , )� ܰ )�  ܰ )�  � )� � )� ܰ +  ,VR_NO_BUS       1    , *~� ܰ *�@ ܰ *�@ � *~� � *~� ܰ +  ,VR_NO_BUS       1    , +:h ܰ +U� ܰ +U� � +:h � +:h ܰ +  ,VR_NO_BUS       1    , ,K� ܰ ,O� ܰ ,O� � ,K� � ,K� ܰ +  ,VR_NO_BUS       1    , - � ܰ -I� ܰ -I� � - � � - � ܰ +  ,VR_NO_BUS       1    , .?� ܰ /�h ܰ /�h � .?� � .?� ܰ +  ,VR_NO_BUS       1    , o0 ܰ Q� ܰ Q� � o0 � o0 ܰ +  ,VR_NO_BUS       1    , "� $� ,� $� ,� K� "� K� "� $� +  ,VR_NO_BUS       1    , @� ܰ J� ܰ J� � @� � @� ܰ +  ,VR_NO_BUS       1    , �h ܰ �� ܰ �� � �h � �h ܰ +  ,VR_NO_BUS       1    , �� ܰ �� ܰ �� � �� � �� ܰ +  ,VR_NO_BUS       1    , #h ܰ >� ܰ >� � #h � #h ܰ +  ,VR_NO_BUS       1    , �( ܰ � ܰ � � �( � �( ܰ +  ,VR_NO_BUS       1    , � ܰ � ܰ � � � � � ܰ +  ,VR_NO_BUS       1    , �h ܰ �� ܰ �� � �h � �h ܰ +  ,VR_NO_BUS       1    , O� ܰ k@ ܰ k@ � O� � O� ܰ +  ,VR_NO_BUS       1    , aX ܰ e@ ܰ e@ � aX � aX ܰ +  ,VR_NO_BUS       1    , 6< ܰ @  ܰ @  � 6< � 6< ܰ +  ,VR_NO_BUS       1    , �� ܰ �@ ܰ �@ � �� � �� ܰ +  ,VR_NO_BUS       1    ,  �X ܰ  �@ ܰ  �@ �  �X �  �X ܰ +  ,VR_NO_BUS       1    , !�< ܰ !�  ܰ !�  � !�< � !�< ܰ +  ,VR_NO_BUS       1    , "1� ܰ "M@ ܰ "M@ � "1� � "1� ܰ +  ,VR_NO_BUS       1    , #CX ܰ #G@ ܰ #G@ � #CX � #CX ܰ +  ,VR_NO_BUS       1    , � ܰ � ܰ � � � � � ܰ +  ,VR_NO_BUS       1    , � ܰ �� ܰ �� � � � � ܰ +  ,VR_NO_BUS       1    , �| ܰ �@ ܰ �@ � �| � �| ܰ +  ,VR_NO_BUS       1    , ,� ܰ H@ ܰ H@ � ,� � ,� ܰ +  ,VR_NO_BUS       1    , �� ܰ �@ ܰ �@ � �� � �� ܰ +  ,VR_NO_BUS       1    , �< ܰ �  ܰ �  � �< � �< ܰ +  ,VR_NO_BUS       1    , p� ܰ z� ܰ z� � p� � p� ܰ +  ,VR_NO_BUS       1    , p� ܰ t� ܰ t� � p� � p� ܰ +  ,VR_NO_BUS       1    , E� ܰ O� ܰ O� � E� � E� ܰ +  ,VR_NO_BUS       1    , E� ܰ I� ܰ I� � E� � E� ܰ +  ,VR_NO_BUS       1    , | ܰ $@ ܰ $@ � | � | ܰ +  ,VR_NO_BUS       1    , X ܰ @ ܰ @ � X � X ܰ +  ,VR_NO_BUS       1    , �< ܰ �  ܰ �  � �< � �< ܰ +  ,VR_NO_BUS       1    , Z� ܰ v  ܰ v  � Z� � Z� ܰ +  ,VR_NO_BUS       1    , l ܰ p  ܰ p  � l � l ܰ +  ,VR_NO_BUS       1    , -� wh -�  wh -�  �x -� �x -� wh +  ,VR_NO_BUS       1    , .f� wh /�h wh /�h �x .f� �x .f� wh +  ,VR_NO_BUS       1    , o0 wh Q� wh Q� �x o0 �x o0 wh +  ,VR_NO_BUS       1    , Ҩ ܰ �  ܰ �  � Ҩ � Ҩ ܰ +  ,VR_NO_BUS       1    , � ܰ �  ܰ �  � � � � ܰ +  ,VR_NO_BUS       1    , �h ܰ �� ܰ �� � �h � �h ܰ +  ,VR_NO_BUS       1    , $h ܰ ?� ܰ ?� � $h � $h ܰ +  ,VR_NO_BUS       1    , �( ܰ � ܰ � � �( � �( ܰ +  ,VR_NO_BUS       1    , � ܰ � ܰ � � � � � ܰ +  ,VR_NO_BUS       1    , �� ܰ �  ܰ �  � �� � �� ܰ +  ,VR_NO_BUS       1    , P� ܰ l@ ܰ l@ � P� � P� ܰ +  ,VR_NO_BUS       1    , 	=< ܰ 	G  ܰ 	G  � 	=< � 	=< ܰ +  ,VR_NO_BUS       1    , 	�� ܰ 	�  ܰ 	�  � 	�� � 	�� ܰ +  ,VR_NO_BUS       1    , 
� ܰ 
�  ܰ 
�  � 
� � 
� ܰ +  ,VR_NO_BUS       1    , � ܰ ;  ܰ ;  � � � � ܰ +  ,VR_NO_BUS       1    ,  �� wh  �@ wh  �@ �x  �� �x  �� wh +  ,VR_NO_BUS       1    , !�X wh !�@ wh !�@ �x !�X �x !�X wh +  ,VR_NO_BUS       1    , "�� wh "�@ wh "�@ �x "�� �x "�� wh +  ,VR_NO_BUS       1    , #+� wh #G@ wh #G@ �x #+� �x #+� wh +  ,VR_NO_BUS       1    , $=X wh $A@ wh $A@ �x $=X �x $=X wh +  ,VR_NO_BUS       1    , $�( wh $݀ wh $݀ �x $�( �x $�( wh +  ,VR_NO_BUS       1    , %�| wh %�@ wh %�@ �x %�| �x %�| wh +  ,VR_NO_BUS       1    , &�< wh &�  wh &�  �x &�< �x &�< wh +  ,VR_NO_BUS       1    , '� wh '�  wh '�  �x '� �x '� wh +  ,VR_NO_BUS       1    , (� wh (�  wh (�  �x (� �x (� wh +  ,VR_NO_BUS       1    , )W� wh )a� wh )a� �x )W� �x )W� wh +  ,VR_NO_BUS       1    , *W� wh *[� wh *[� �x *W� �x *W� wh +  ,VR_NO_BUS       1    , +Q� wh +�@ wh +�@ �x +Q� �x +Q� wh +  ,VR_NO_BUS       1    , ,4h wh ,O� wh ,O� �x ,4h �x ,4h wh +  ,VR_NO_BUS       1    , ,Ш wh ,�  wh ,�  �x ,Ш �x ,Ш wh +  ,VR_NO_BUS       1    , �( wh ƀ wh ƀ �x �( �x �( wh +  ,VR_NO_BUS       1    , �� wh �� wh �� �x �� �x �� wh +  ,VR_NO_BUS       1    , �| wh �@ wh �@ �x �| �x �| wh +  ,VR_NO_BUS       1    , l< wh v  wh v  �x l< �x l< wh +  ,VR_NO_BUS       1    , ר wh �  wh �  �x ר �x ר wh +  ,VR_NO_BUS       1    , � wh �  wh �  �x � �x � wh +  ,VR_NO_BUS       1    , �� wh �� wh �� �x �� �x �� wh +  ,VR_NO_BUS       1    , �� wh �� wh �� �x �� �x �� wh +  ,VR_NO_BUS       1    , �� wh �� wh �� �x �� �x �� wh +  ,VR_NO_BUS       1    , �� wh �� wh �� �x �� �x �� wh +  ,VR_NO_BUS       1    , �� wh �� wh �� �x �� �x �� wh +  ,VR_NO_BUS       1    , a| wh k@ wh k@ �x a| �x a| wh +  ,VR_NO_BUS       1    , aX wh e@ wh e@ �x aX �x aX wh +  ,VR_NO_BUS       1    , [X wh _@ wh _@ �x [X �x [X wh +  ,VR_NO_BUS       1    , �h wh  � wh  � �x �h �x �h wh +  ,VR_NO_BUS       1    , 
� wh � wh � �x 
� �x 
� wh +  ,VR_NO_BUS       1    , 
� wh � wh � �x 
� �x 
� wh +  ,VR_NO_BUS       1    , �h wh �� wh �� �x �h �x �h wh +  ,VR_NO_BUS       1    , 	�\ wh 	�� wh 	�� �x 	�\ �x 	�\ wh +  ,VR_NO_BUS       1    , 
�\ wh 
�� wh 
�� �x 
�\ �x 
�\ wh +  ,VR_NO_BUS       1    , o� wh y� wh y� �x o� �x o� wh +  ,VR_NO_BUS       1    , �( wh �� wh �� �x �( �x �( wh +  ,VR_NO_BUS       1    , �| wh �@ wh �@ �x �| �x �| wh +  ,VR_NO_BUS       1    , T wh m� wh m� �x T �x T wh +  ,VR_NO_BUS       1    , �\ wh 	� wh 	� �x �\ �x �\ wh +  ,VR_NO_BUS       1    , ڼ wh � wh � �x ڼ �x ڼ wh +  ,VR_NO_BUS       1    , �h wh �� wh �� �x �h �x �h wh +  ,VR_NO_BUS       1    , �\ wh �� wh �� �x �\ �x �\ wh +  ,VR_NO_BUS       1    , �� wh �@ wh �@ �x �� �x �� wh +  ,VR_NO_BUS       1    , �� wh �@ wh �@ �x �� �x �� wh +  ,VR_NO_BUS       1    , &�( 
L� &р 
L� &р 
s� &�( 
s� &�( 
L� +  ,VR_NO_BUS       1    , 'ǘ 
L� 'ˀ 
L� 'ˀ 
s� 'ǘ 
s� 'ǘ 
L� +  ,VR_NO_BUS       1    , (�| 
L� (�@ 
L� (�@ 
s� (�| 
s� (�| 
L� +  ,VR_NO_BUS       1    , )w< 
L� )�  
L� )�  
s� )w< 
s� )w< 
L� +  ,VR_NO_BUS       1    , *w 
L� *{  
L� *{  
s� *w 
s� *w 
L� +  ,VR_NO_BUS       1    , +q 
L� +u  
L� +u  
s� +q 
s� +q 
L� +  ,VR_NO_BUS       1    , ,k 
L� ,o  
L� ,o  
s� ,k 
s� ,k 
L� +  ,VR_NO_BUS       1    , -e 
L� -i  
L� -i  
s� -e 
s� -e 
L� +  ,VR_NO_BUS       1    , .9� 
L� /�h 
L� /�h 
s� .9� 
s� .9� 
L� +  ,VR_NO_BUS       1    , o0 
L� Q� 
L� Q� 
s� o0 
s� o0 
L� +  ,VR_NO_BUS       1    , G� wh K� wh K� �x G� �x G� wh +  ,VR_NO_BUS       1    , �� wh @ wh @ �x �� �x �� wh +  ,VR_NO_BUS       1    , �( wh �� wh �� �x �( �x �( wh +  ,VR_NO_BUS       1    , �� wh �� wh �� �x �� �x �� wh +  ,VR_NO_BUS       1    , h wh 9� wh 9� �x h �x h wh +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , m| 
L� w@ 
L� w@ 
s� m| 
s� m| 
L� +  ,VR_NO_BUS       1    , H< 
L� R  
L� R  
s� H< 
s� H< 
L� +  ,VR_NO_BUS       1    , "� 
L� ,� 
L� ,� 
s� "� 
s� "� 
L� +  ,VR_NO_BUS       1    , "� 
L� &� 
L� &� 
s� "� 
s� "� 
L� +  ,VR_NO_BUS       1    , �� 
L� �@ 
L� �@ 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , �h 
L� �� 
L� �� 
s� �h 
s� �h 
L� +  ,VR_NO_BUS       1    ,  n� 
L�  x� 
L�  x� 
s�  n� 
s�  n� 
L� +  ,VR_NO_BUS       1    , !n� 
L� !r� 
L� !r� 
s� !n� 
s� !n� 
L� +  ,VR_NO_BUS       1    , "C| 
L� "M@ 
L� "M@ 
s� "C| 
s� "C| 
L� +  ,VR_NO_BUS       1    , #CX 
L� #G@ 
L� #G@ 
s� #CX 
s� #CX 
L� +  ,VR_NO_BUS       1    , #�� 
L� #�@ 
L� #�@ 
s� #�� 
s� #�� 
L� +  ,VR_NO_BUS       1    , $�X 
L� $�@ 
L� $�@ 
s� $�X 
s� $�X 
L� +  ,VR_NO_BUS       1    , %}� 
L� %�  
L� %�  
s� %}� 
s� %}� 
L� +  ,VR_NO_BUS       1    , &9( 
L� &T� 
L� &T� 
s� &9( 
s� &9( 
L� +  ,VR_NO_BUS       1    , �( 
L� � 
L� � 
s� �( 
s� �( 
L� +  ,VR_NO_BUS       1    , �� 
L� �@ 
L� �@ 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    ,  � 
L� <@ 
L� <@ 
s�  � 
s�  � 
L� +  ,VR_NO_BUS       1    , < 
L�   
L�   
s� < 
s� < 
L� +  ,VR_NO_BUS       1    , x� 
L� �  
L� �  
s� x� 
s� x� 
L� +  ,VR_NO_BUS       1    , �� 
L�   
L�   
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , � 
L� ̀ 
L� ̀ 
s� � 
s� � 
L� +  ,VR_NO_BUS       1    , �| 
L� �@ 
L� �@ 
s� �| 
s� �| 
L� +  ,VR_NO_BUS       1    , � 
L� $@ 
L� $@ 
s� � 
s� � 
L� +  ,VR_NO_BUS       1    , � 
L� @ 
L� @ 
s� � 
s� � 
L� +  ,VR_NO_BUS       1    , �< 
L� �  
L� �  
s� �< 
s� �< 
L� +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , o0 " Q� " Q� I o0 I o0 " +  ,VR_NO_BUS       1    , Ҩ 
L� �  
L� �  
s� Ҩ 
s� Ҩ 
L� +  ,VR_NO_BUS       1    , � 
L� �  
L� �  
s� � 
s� � 
L� +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , �� 
L� �� 
L� �� 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , b| 
L� l@ 
L� l@ 
s� b| 
s� b| 
L� +  ,VR_NO_BUS       1    , 	=< 
L� 	G  
L� 	G  
s� 	=< 
s� 	=< 
L� +  ,VR_NO_BUS       1    , 
D� 
L� 
`@ 
L� 
`@ 
s� 
D� 
s� 
D� 
L� +  ,VR_NO_BUS       1    , 
�� 
L� 
�@ 
L� 
�@ 
s� 
�� 
s� 
�� 
L� +  ,VR_NO_BUS       1    , �( 
L� �� 
L� �� 
s� �( 
s� �( 
L� +  ,VR_NO_BUS       1    , �� 
L� �@ 
L� �@ 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , 2� 
L� N@ 
L� N@ 
s� 2� 
s� 2� 
L� +  ,VR_NO_BUS       1    , �� 
L� �@ 
L� �@ 
s� �� 
s� �� 
L� +  ,VR_NO_BUS       1    , !� " !� " !� I !� I !� " +  ,VR_NO_BUS       1    , "�| " "�@ " "�@ I "�| I "�| " +  ,VR_NO_BUS       1    , #�X " #�@ " #�@ I #�X I #�X " +  ,VR_NO_BUS       1    , $�X " $�@ " $�@ I $�X I $�X " +  ,VR_NO_BUS       1    , %�X " %�@ " %�@ I %�X I %�X " +  ,VR_NO_BUS       1    , &w� " &�  " &�  I &w� I &w� " +  ,VR_NO_BUS       1    , '� " '�  " '�  I '� I '� " +  ,VR_NO_BUS       1    , (]� " (g� " (g� I (]� I (]� " +  ,VR_NO_BUS       1    , )]� " )a� " )a� I )]� I )]� " +  ,VR_NO_BUS       1    , )� " )�  " )�  I )� I )� " +  ,VR_NO_BUS       1    , *�� " *�� " *�� I *�� I *�� " +  ,VR_NO_BUS       1    , +�� " +�� " +�� I +�� I +�� " +  ,VR_NO_BUS       1    , ,�� " ,�� " ,�� I ,�� I ,�� " +  ,VR_NO_BUS       1    , -~| " -�@ " -�@ I -~| I -~| " +  ,VR_NO_BUS       1    , .~X " /�h " /�h I .~X I .~X " +  ,VR_NO_BUS       1    , �( " �� " �� I �( I �( " +  ,VR_NO_BUS       1    , �h " �� " �� I �h I �h " +  ,VR_NO_BUS       1    , �( " �� " �� I �( I �( " +  ,VR_NO_BUS       1    , �h " �� " �� I �h I �h " +  ,VR_NO_BUS       1    , /h " J� " J� I /h I /h " +  ,VR_NO_BUS       1    , � " %� " %� I � I � " +  ,VR_NO_BUS       1    , �| "  @ "  @ I �| I �| " +  ,VR_NO_BUS       1    , �< " �  " �  I �< I �< " +  ,VR_NO_BUS       1    , � " �  " �  I � I � " +  ,VR_NO_BUS       1    , � " �  " �  I � I � " +  ,VR_NO_BUS       1    , �� " �� " �� I �� I �� " +  ,VR_NO_BUS       1    , *� " F  " F  I *� I *� " +  ,VR_NO_BUS       1    , � "  � "  � I � I � " +  ,VR_NO_BUS       1    ,  � "  � "  � I  � I  � " +  ,VR_NO_BUS       1    ,  � "  �� "  �� I  � I  � " +  ,VR_NO_BUS       1    , 
�� " 
�  " 
�  I 
�� I 
�� " +  ,VR_NO_BUS       1    , ^( " y� " y� I ^( I ^( " +  ,VR_NO_BUS       1    , �( " �� " �� I �( I �( " +  ,VR_NO_BUS       1    , �| " �@ " �@ I �| I �| " +  ,VR_NO_BUS       1    , �< " �  " �  I �< I �< " +  ,VR_NO_BUS       1    , � " �  " �  I � I � " +  ,VR_NO_BUS       1    , � " #  " #  I � I � " +  ,VR_NO_BUS       1    , �� " �@ " �@ I �� I �� " +  ,VR_NO_BUS       1    ,  � " <@ " <@ I  � I  � " +  ,VR_NO_BUS       1    , �( " ؀ " ؀ I �( I �( " +  ,VR_NO_BUS       1    , :( " U� " U� I :( I :( " +  ,VR_NO_BUS       1    , �( " Ҁ " Ҁ I �( I �( " +  ,VR_NO_BUS       1    , 4( " O� " O� I 4( I 4( " +  ,VR_NO_BUS       1    , � " *@ " *@ I � I � " +  ,VR_NO_BUS       1    , (( " C� " C� I (( I (( " +  ,VR_NO_BUS       1    , *_� � *{  � *{  A� *_� A� *_� � +  ,VR_NO_BUS       1    , *�� � +@ � +@ A� *�� A� *�� � +  ,VR_NO_BUS       1    , +�h � +�� � +�� A� +�h A� +�h � +  ,VR_NO_BUS       1    , ,r� � ,�@ � ,�@ A� ,r� A� ,r� � +  ,VR_NO_BUS       1    , -.h � /�h � /�h A� -.h A� -.h � +  ,VR_NO_BUS       1    , o0 � Q� � Q� A� o0 A� o0 � +  ,VR_NO_BUS       1    , Ҩ " �  " �  I Ҩ I Ҩ " +  ,VR_NO_BUS       1    , �� " �� " �� I �� I �� " +  ,VR_NO_BUS       1    , �� " �� " �� I �� I �� " +  ,VR_NO_BUS       1    , �� " �� " �� I �� I �� " +  ,VR_NO_BUS       1    , n| " x@ " x@ I n| I n| " +  ,VR_NO_BUS       1    , I< " S  " S  I I< I I< " +  ,VR_NO_BUS       1    , �� " �  " �  I �� I �� " +  ,VR_NO_BUS       1    , �� " �� " �� I �� I �� " +  ,VR_NO_BUS       1    , 	�� " 	�� " 	�� I 	�� I 	�� " +  ,VR_NO_BUS       1    , "� � &� � &� A� "� A� "� � +  ,VR_NO_BUS       1    , � �  � �  � A� � A� � � +  ,VR_NO_BUS       1    , � � �� � �� A� � A� � � +  ,VR_NO_BUS       1    ,  � �  �� �  �� A�  � A�  � � +  ,VR_NO_BUS       1    , !� � !� � !� A� !� A� !� � +  ,VR_NO_BUS       1    , "�| � "�@ � "�@ A� "�| A� "�| � +  ,VR_NO_BUS       1    , #�< � #�  � #�  A� #�< A� #�< � +  ,VR_NO_BUS       1    , $%� � $A@ � $A@ A� $%� A� $%� � +  ,VR_NO_BUS       1    , $�� � $�@ � $�@ A� $�� A� $�� � +  ,VR_NO_BUS       1    , %�X � %�@ � %�@ A� %�X A� %�X � +  ,VR_NO_BUS       1    , &9( � &T� � &T� A� &9( A� &9( � +  ,VR_NO_BUS       1    , '%| � '/@ � '/@ A� '%| A� '%| � +  ,VR_NO_BUS       1    , (%X � ()@ � ()@ A� (%X A� (%X � +  ,VR_NO_BUS       1    , )X � )#@ � )#@ A� )X A� )X � +  ,VR_NO_BUS       1    , )�( � )�� � )�� A� )�( A� )�( � +  ,VR_NO_BUS       1    , �� � �@ � �@ A� �� A� �� � +  ,VR_NO_BUS       1    , �X � �@ � �@ A� �X A� �X � +  ,VR_NO_BUS       1    , ~< � �  � �  A� ~< A� ~< � +  ,VR_NO_BUS       1    , ~ � �  � �  A� ~ A� ~ � +  ,VR_NO_BUS       1    , R� � \� � \� A� R� A� R� � +  ,VR_NO_BUS       1    , R� � V� � V� A� R� A� R� � +  ,VR_NO_BUS       1    , L� � P� � P� A� L� A� L� � +  ,VR_NO_BUS       1    , �h � �� � �� A� �h A� �h � +  ,VR_NO_BUS       1    , �� � �� � �� A� �� A� �� � +  ,VR_NO_BUS       1    , �� � �� � �� A� �� A� �� � +  ,VR_NO_BUS       1    , B� � ^  � ^  A� B� A� B� � +  ,VR_NO_BUS       1    , .� � 8� � 8� A� .� A� .� � +  ,VR_NO_BUS       1    , �h � �� � �� A� �h A� �h � +  ,VR_NO_BUS       1    , 6� � R  � R  A� 6� A� 6� � +  ,VR_NO_BUS       1    , "� � ,� � ,� A� "� A� "� � +  ,VR_NO_BUS       1    , �( � �� � �� A� �( A� �( � +  ,VR_NO_BUS       1    , n| � x@ � x@ A� n| A� n| � +  ,VR_NO_BUS       1    , nX � r@ � r@ A� nX A� nX � +  ,VR_NO_BUS       1    , C< � M  � M  A� C< A� C< � +  ,VR_NO_BUS       1    , 	� � 	'� � 	'� A� 	� A� 	� � +  ,VR_NO_BUS       1    , 
� � 
!� � 
!� A� 
� A� 
� � +  ,VR_NO_BUS       1    , 
�h � 
�� � 
�� A� 
�h A� 
�h � +  ,VR_NO_BUS       1    ,  h � � � � A�  h A�  h � +  ,VR_NO_BUS       1    , � � �� � �� A� � A� � � +  ,VR_NO_BUS       1    , � � �� � �� A� � A� � � +  ,VR_NO_BUS       1    , �| � �@ � �@ A� �| A� �| � +  ,VR_NO_BUS       1    , �< � �  � �  A� �< A� �< � +  ,VR_NO_BUS       1    , � � �  � �  A� � A� � � +  ,VR_NO_BUS       1    , p� � z� � z� A� p� A� p� � +  ,VR_NO_BUS       1    , � � 6@ � 6@ A� � A� � � +  ,VR_NO_BUS       1    , #�h А $� А $� �� #�h �� #�h А +  ,VR_NO_BUS       1    , $dh А $� А $� �� $dh �� $dh А +  ,VR_NO_BUS       1    , %u� А %y� А %y� �� %u� �� %u� А +  ,VR_NO_BUS       1    , &� А &5@ А &5@ �� &� �� &� А +  ,VR_NO_BUS       1    , '+X А '/@ А '/@ �� '+X �� '+X А +  ,VR_NO_BUS       1    , ( < А (
  А (
  �� ( < �� ( < А +  ,VR_NO_BUS       1    , )  А )  А )  �� )  �� )  А +  ,VR_NO_BUS       1    , )�� А )�@ А )�@ �� )�� �� )�� А +  ,VR_NO_BUS       1    , *@h А *[� А *[� �� *@h �� *@h А +  ,VR_NO_BUS       1    , *�� А +@ А +@ �� *�� �� *�� А +  ,VR_NO_BUS       1    , ,X А /�h А /�h �� ,X �� ,X А +  ,VR_NO_BUS       1    , o0 А Q� А Q� �� o0 �� o0 А +  ,VR_NO_BUS       1    , G� � K� � K� A� G� A� G� � +  ,VR_NO_BUS       1    , A� � E� � E� A� A� A� A� � +  ,VR_NO_BUS       1    , ( �  � �  � A� ( A� ( � +  ,VR_NO_BUS       1    , �� А �� А �� �� �� �� �� А +  ,VR_NO_BUS       1    , �� А �� А �� �� �� �� �� А +  ,VR_NO_BUS       1    , /h А J� А J� �� /h �� /h А +  ,VR_NO_BUS       1    , � А %� А %� �� � �� � А +  ,VR_NO_BUS       1    , �| А  @ А  @ �� �| �� �| А +  ,VR_NO_BUS       1    , �< А �  А �  �� �< �� �< А +  ,VR_NO_BUS       1    , � А �  А �  �� � �� � А +  ,VR_NO_BUS       1    , �� А �� А �� �� �� �� �� А +  ,VR_NO_BUS       1    , �� А �� А �� �� �� �� �� А +  ,VR_NO_BUS       1    , z� А �� А �� �� z� �� z� А +  ,VR_NO_BUS       1    , U| А _@ А _@ �� U| �� U| А +  ,VR_NO_BUS       1    ,  UX А  Y@ А  Y@ ��  UX ��  UX А +  ,VR_NO_BUS       1    , !*< А !4  А !4  �� !*< �� !*< А +  ,VR_NO_BUS       1    , "* А ".  А ".  �� "* �� "* А +  ,VR_NO_BUS       1    , #$ А #(  А #(  �� #$ �� #$ А +  ,VR_NO_BUS       1    , 
� А 
�  А 
�  �� 
� �� 
� А +  ,VR_NO_BUS       1    , �� А �� А �� �� �� �� �� А +  ,VR_NO_BUS       1    , �h А � А � �� �h �� �h А +  ,VR_NO_BUS       1    , � А � А � �� � �� � А +  ,VR_NO_BUS       1    , � А 	� А 	� �� � �� � А +  ,VR_NO_BUS       1    , kh А �� А �� �� kh �� kh А +  ,VR_NO_BUS       1    , W� А a� А a� �� W� �� W� А +  ,VR_NO_BUS       1    , 2| А <@ А <@ �� 2| �� 2| А +  ,VR_NO_BUS       1    , 2X А 6@ А 6@ �� 2X �� 2X А +  ,VR_NO_BUS       1    , < А   А   �� < �� < А +  ,VR_NO_BUS       1    , r� А �  А �  �� r� �� r� А +  ,VR_NO_BUS       1    , � А �  А �  �� � �� � А +  ,VR_NO_BUS       1    , X� А b� А b� �� X� �� X� А +  ,VR_NO_BUS       1    , 3� А =� А =� �� 3� �� 3� А +  ,VR_NO_BUS       1    , �( А �� А �� �� �( �� �( А +  ,VR_NO_BUS       1    , '�� � '�� � '�� � '�� � '�� � +  ,VR_NO_BUS       1    , (�� � (ŀ � (ŀ � (�� � (�� � +  ,VR_NO_BUS       1    , )�� � )�� � )�� � )�� � )�� � +  ,VR_NO_BUS       1    , *_� � *{  � *{  � *_� � *_� � +  ,VR_NO_BUS       1    , +( � /�h � /�h � +( � +( � +  ,VR_NO_BUS       1    , o0 � Q� � Q� � o0 � o0 � +  ,VR_NO_BUS       1    , G� А K� А K� �� G� �� G� А +  ,VR_NO_BUS       1    , ( А &� А &� �� ( �� ( А +  ,VR_NO_BUS       1    , �( А �� А �� �� �( �� �( А +  ,VR_NO_BUS       1    , �� А �� А �� �� �� �� �� А +  ,VR_NO_BUS       1    , n| А x@ А x@ �� n| �� n| А +  ,VR_NO_BUS       1    , nX А r@ А r@ �� nX �� nX А +  ,VR_NO_BUS       1    , �� А �@ А �@ �� �� �� �� А +  ,VR_NO_BUS       1    , �X А �@ А �@ �� �X �� �X А +  ,VR_NO_BUS       1    , 	�< А 	�  А 	�  �� 	�< �� 	�< А +  ,VR_NO_BUS       1    , s| � }@ � }@ � s| � s| � +  ,VR_NO_BUS       1    , sX � w@ � w@ � sX � sX � +  ,VR_NO_BUS       1    , H< � R  � R  � H< � H< � +  ,VR_NO_BUS       1    , "� � ,� � ,� � "� � "� � +  ,VR_NO_BUS       1    , �� � � � � � �� � �� � +  ,VR_NO_BUS       1    , �� � � � � � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    ,  �| �  �@ �  �@ �  �| �  �| � +  ,VR_NO_BUS       1    , !�X � !�@ � !�@ � !�X � !�X � +  ,VR_NO_BUS       1    , "�< � "�  � "�  � "�< � "�< � +  ,VR_NO_BUS       1    , #� � #�  � #�  � #� � #� � +  ,VR_NO_BUS       1    , $u� � $� � $� � $u� � $u� � +  ,VR_NO_BUS       1    , %u� � %y� � %y� � %u� � %u� � +  ,VR_NO_BUS       1    , &o� � &s� � &s� � &o� � &o� � +  ,VR_NO_BUS       1    , &�� � '  � '  � &�� � &�� � +  ,VR_NO_BUS       1    , � � �� � �� � � � � � +  ,VR_NO_BUS       1    , � � � � � � � � � � +  ,VR_NO_BUS       1    , �| � �@ � �@ � �| � �| � +  ,VR_NO_BUS       1    , �< � �  � �  � �< � �< � +  ,VR_NO_BUS       1    , � � �  � �  � � � � � +  ,VR_NO_BUS       1    , j� � t� � t� � j� � j� � +  ,VR_NO_BUS       1    , E� � O� � O� � E� � E� � +  ,VR_NO_BUS       1    , E� � I� � I� � E� � E� � +  ,VR_NO_BUS       1    , | � $@ � $@ � | � | � +  ,VR_NO_BUS       1    , X � @ � @ � X � X � +  ,VR_NO_BUS       1    , �< � �  � �  � �< � �< � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , �� � �� � �� � �� � �� � +  ,VR_NO_BUS       1    , `� "�\  "�\  "� `� "� `� "�\      1    , �� �� � �� � �� �� �� �� ��      1    , � � � � � �� � �� � �      1    , G� � K� � K� � G� � G� � +  ,VR_NO_BUS       1    , �h � �� � �� � �h � �h � +  ,VR_NO_BUS       1    , �( � �� � �� � �( � �( � +  ,VR_NO_BUS       1    , ( �  � �  � � ( � ( � +  ,VR_NO_BUS       1    , � � � � � � � � � � +  ,VR_NO_BUS       1    , �| � �@ � �@ � �| � �| � +  ,VR_NO_BUS       1    , �X � �@ � �@ � �X � �X � +  ,VR_NO_BUS       1    , �� � �  � �  � �� � �� � +  ,VR_NO_BUS       1    , 	+� � 	G  � 	G  � 	+� � 	+� � +  ,VR_NO_BUS       1    , 
� � 
!� � 
!� � 
� � 
� � +  ,VR_NO_BUS       1    , � � � � � � � � � � +  ,VR_NO_BUS       1    , �( � �� � �� � �( � �( � +  ,VR_NO_BUS       
       $�L &�x 
CLOCK       
       %+� &�x 
RESET              0� #۰ I_VALID              0� $� 
READY       
       #EL &�x O_VALID               | �� EDGE              | � VDD       
       *�\  	� 
T22[0]             0� ' 
T21[1]             0� o 
T21[2]             0� �X 
T22[1]              | �� 
T22[7]              | T` 
T22[6]              | �x 
T21[7]      
       N� &�x 
T22[5]      
       
� &�x 
T21[6]             0� � 
T22[4]      
       �� &�x 
T21[5]             0� �� 
T22[3]             0� 9P 
T21[4]      
       &ɰ  	� 
T22[2]             0� @ 
T21[3]      
       .*\  	� 
T02[0]      
       *B\  	� 
T20[0]      
        ~\  	� 
T21[0]      
       $�  	� 
T20[1]      
       $^�  	� 
T20[2]              | "�� 
T20[7]      
       >� &�x 
T20[6]      
       { &�x 
T20[5]             0�  � 
T20[4]      
       %��  	� 
T20[3]      
        8  	� 
T12[0]      
       &;  	� 
T10[0]      
       ('L  	� 
T10[1]             0� ?� 
T10[2]      
       k� &�x 
T10[7]              | &0 
T10[6]      
       �T &�x 
T10[5]      
       #x &�x 
T10[4]             0� {p 
T10[3]      
       )��  	� 
T00[0]             0� ɔ 
T02[1]             0� � 
T02[2]             0� � 
T12[1]              | �h 
T12[7]              | ܈ 
T02[7]      
       �( &�x 
T12[6]      
       �� &�x 
T02[6]      
       A� &�x 
T12[5]      
       , &�x 
T02[5]             0� T` 
T12[4]             0� � 
T02[4]             0� �( 
T12[3]             0� �X 
T02[3]             0� -P 
T12[2]      
       )�4  	� 
T01[0]      
       �$  	� 
T00[1]             0� �� 
T00[2]      
       	�� &�x 
T00[6]              | %�8 
T00[7]      
       	J� &�x 
T00[5]             0� ؠ 
T00[4]      
       �� &�x 
T00[3]      
       -d  	� 
T01[1]      
       -n�  	� 
T01[2]              | !�8 
T01[7]      
       N� &�x 
T01[6]      
        j� &�x 
T01[5]             0� �� 
T01[4]      
       .UT  	� 
T01[3]             0� � GND               | j� DIRECTION[1]              | ct DIRECTION[0]      
       
�|  	� DIRECTION[2]              | �, THRESHOLD[10]               | #$ THRESHOLD[9]              | =� THRESHOLD[8]              | �� THRESHOLD[7]      
       L  	� THRESHOLD[6]      
       \�  	� THRESHOLD[5]      
       XL  	� THRESHOLD[4]              | �� THRESHOLD[3]              | �� THRESHOLD[2]      
       �� &�x THRESHOLD[1]      
       �� &�x THRESHOLD[0]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              